module result_buffer (
	input CLK,
	input RSTN,
	input i_result_in_en,
	input i_result_out_en,
	input [7:0] i_counter,
	input [31:0] i_data0,
	input [31:0] i_data1,
	input [31:0] i_data2,
	input [31:0] i_data3,
	input [31:0] i_data4,
	input [31:0] i_data5,
	input [31:0] i_data6,
	input [31:0] i_data7,
	input [31:0] i_data8,
	input [31:0] i_data9,
	input [31:0] i_data10,
	input [31:0] i_data11,
	input [31:0] i_data12,
	input [31:0] i_data13,
	input [31:0] i_data14,
	input [31:0] i_data15,
	input [31:0] i_data16,
	input [31:0] i_data17,
	input [31:0] i_data18,
	input [31:0] i_data19,
	input [31:0] i_data20,
	input [31:0] i_data21,
	input [31:0] i_data22,
	input [31:0] i_data23,
	input [31:0] i_data24,
	input [31:0] i_data25,
	input [31:0] i_data26,
	input [31:0] i_data27,
	input [31:0] i_data28,
	input [31:0] i_data29,
	input [31:0] i_data30,
	input [31:0] i_data31,
	input [31:0] i_data32,
	input [31:0] i_data33,
	input [31:0] i_data34,
	input [31:0] i_data35,
	input [31:0] i_data36,
	input [31:0] i_data37,
	input [31:0] i_data38,
	input [31:0] i_data39,
	input [31:0] i_data40,
	input [31:0] i_data41,
	input [31:0] i_data42,
	input [31:0] i_data43,
	input [31:0] i_data44,
	input [31:0] i_data45,
	input [31:0] i_data46,
	input [31:0] i_data47,
	input [31:0] i_data48,
	input [31:0] i_data49,
	input [31:0] i_data50,
	input [31:0] i_data51,
	input [31:0] i_data52,
	input [31:0] i_data53,
	input [31:0] i_data54,
	input [31:0] i_data55,
	input [31:0] i_data56,
	input [31:0] i_data57,
	input [31:0] i_data58,
	input [31:0] i_data59,
	input [31:0] i_data60,
	input [31:0] i_data61,
	input [31:0] i_data62,
	input [31:0] i_data63,
	input [31:0] i_data64,
	input [31:0] i_data65,
	input [31:0] i_data66,
	input [31:0] i_data67,
	input [31:0] i_data68,
	input [31:0] i_data69,
	input [31:0] i_data70,
	input [31:0] i_data71,
	input [31:0] i_data72,
	input [31:0] i_data73,
	input [31:0] i_data74,
	input [31:0] i_data75,
	input [31:0] i_data76,
	input [31:0] i_data77,
	input [31:0] i_data78,
	input [31:0] i_data79,
	input [31:0] i_data80,
	input [31:0] i_data81,
	input [31:0] i_data82,
	input [31:0] i_data83,
	input [31:0] i_data84,
	input [31:0] i_data85,
	input [31:0] i_data86,
	input [31:0] i_data87,
	input [31:0] i_data88,
	input [31:0] i_data89,
	input [31:0] i_data90,
	input [31:0] i_data91,
	input [31:0] i_data92,
	input [31:0] i_data93,
	input [31:0] i_data94,
	input [31:0] i_data95,
	input [31:0] i_data96,
	input [31:0] i_data97,
	input [31:0] i_data98,
	input [31:0] i_data99,
	input [31:0] i_data100,
	input [31:0] i_data101,
	input [31:0] i_data102,
	input [31:0] i_data103,
	input [31:0] i_data104,
	input [31:0] i_data105,
	input [31:0] i_data106,
	input [31:0] i_data107,
	input [31:0] i_data108,
	input [31:0] i_data109,
	input [31:0] i_data110,
	input [31:0] i_data111,
	input [31:0] i_data112,
	input [31:0] i_data113,
	input [31:0] i_data114,
	input [31:0] i_data115,
	input [31:0] i_data116,
	input [31:0] i_data117,
	input [31:0] i_data118,
	input [31:0] i_data119,
	input [31:0] i_data120,
	input [31:0] i_data121,
	input [31:0] i_data122,
	input [31:0] i_data123,
	input [31:0] i_data124,
	input [31:0] i_data125,
	input [31:0] i_data126,
	input [31:0] i_data127,
	input [31:0] i_data128,
	input [31:0] i_data129,
	input [31:0] i_data130,
	input [31:0] i_data131,
	input [31:0] i_data132,
	input [31:0] i_data133,
	input [31:0] i_data134,
	input [31:0] i_data135,
	input [31:0] i_data136,
	input [31:0] i_data137,
	input [31:0] i_data138,
	input [31:0] i_data139,
	input [31:0] i_data140,
	input [31:0] i_data141,
	input [31:0] i_data142,
	input [31:0] i_data143,
	input [31:0] i_data144,
	input [31:0] i_data145,
	input [31:0] i_data146,
	input [31:0] i_data147,
	input [31:0] i_data148,
	input [31:0] i_data149,
	input [31:0] i_data150,
	input [31:0] i_data151,
	input [31:0] i_data152,
	input [31:0] i_data153,
	input [31:0] i_data154,
	input [31:0] i_data155,
	input [31:0] i_data156,
	input [31:0] i_data157,
	input [31:0] i_data158,
	input [31:0] i_data159,
	input [31:0] i_data160,
	input [31:0] i_data161,
	input [31:0] i_data162,
	input [31:0] i_data163,
	input [31:0] i_data164,
	input [31:0] i_data165,
	input [31:0] i_data166,
	input [31:0] i_data167,
	input [31:0] i_data168,
	input [31:0] i_data169,
	input [31:0] i_data170,
	input [31:0] i_data171,
	input [31:0] i_data172,
	input [31:0] i_data173,
	input [31:0] i_data174,
	input [31:0] i_data175,
	input [31:0] i_data176,
	input [31:0] i_data177,
	input [31:0] i_data178,
	input [31:0] i_data179,
	input [31:0] i_data180,
	input [31:0] i_data181,
	input [31:0] i_data182,
	input [31:0] i_data183,
	input [31:0] i_data184,
	input [31:0] i_data185,
	input [31:0] i_data186,
	input [31:0] i_data187,
	input [31:0] i_data188,
	input [31:0] i_data189,
	input [31:0] i_data190,
	input [31:0] i_data191,
	input [31:0] i_data192,
	input [31:0] i_data193,
	input [31:0] i_data194,
	input [31:0] i_data195,
	input [31:0] i_data196,
	input [31:0] i_data197,
	input [31:0] i_data198,
	input [31:0] i_data199,
	input [31:0] i_data200,
	input [31:0] i_data201,
	input [31:0] i_data202,
	input [31:0] i_data203,
	input [31:0] i_data204,
	input [31:0] i_data205,
	input [31:0] i_data206,
	input [31:0] i_data207,
	input [31:0] i_data208,
	input [31:0] i_data209,
	input [31:0] i_data210,
	input [31:0] i_data211,
	input [31:0] i_data212,
	input [31:0] i_data213,
	input [31:0] i_data214,
	input [31:0] i_data215,
	input [31:0] i_data216,
	input [31:0] i_data217,
	input [31:0] i_data218,
	input [31:0] i_data219,
	input [31:0] i_data220,
	input [31:0] i_data221,
	input [31:0] i_data222,
	input [31:0] i_data223,
	input [31:0] i_data224,
	input [31:0] i_data225,
	input [31:0] i_data226,
	input [31:0] i_data227,
	input [31:0] i_data228,
	input [31:0] i_data229,
	input [31:0] i_data230,
	input [31:0] i_data231,
	input [31:0] i_data232,
	input [31:0] i_data233,
	input [31:0] i_data234,
	input [31:0] i_data235,
	input [31:0] i_data236,
	input [31:0] i_data237,
	input [31:0] i_data238,
	input [31:0] i_data239,
	input [31:0] i_data240,
	input [31:0] i_data241,
	input [31:0] i_data242,
	input [31:0] i_data243,
	input [31:0] i_data244,
	input [31:0] i_data245,
	input [31:0] i_data246,
	input [31:0] i_data247,
	input [31:0] i_data248,
	input [31:0] i_data249,
	input [31:0] i_data250,
	input [31:0] i_data251,
	input [31:0] i_data252,
	input [31:0] i_data253,
	input [31:0] i_data254,
	input [31:0] i_data255,
	output [31:0] o_data
);

	reg [31:0] buffer [0:255];

	always @(posedge CLK) begin
		if (!RSTN) begin
			buffer[  0] <= 0;
			buffer[  1] <= 0;
			buffer[  2] <= 0;
			buffer[  3] <= 0;
			buffer[  4] <= 0;
			buffer[  5] <= 0;
			buffer[  6] <= 0;
			buffer[  7] <= 0;
			buffer[  8] <= 0;
			buffer[  9] <= 0;
			buffer[ 10] <= 0;
			buffer[ 11] <= 0;
			buffer[ 12] <= 0;
			buffer[ 13] <= 0;
			buffer[ 14] <= 0;
			buffer[ 15] <= 0;
			buffer[ 16] <= 0;
			buffer[ 17] <= 0;
			buffer[ 18] <= 0;
			buffer[ 19] <= 0;
			buffer[ 20] <= 0;
			buffer[ 21] <= 0;
			buffer[ 22] <= 0;
			buffer[ 23] <= 0;
			buffer[ 24] <= 0;
			buffer[ 25] <= 0;
			buffer[ 26] <= 0;
			buffer[ 27] <= 0;
			buffer[ 28] <= 0;
			buffer[ 29] <= 0;
			buffer[ 30] <= 0;
			buffer[ 31] <= 0;
			buffer[ 32] <= 0;
			buffer[ 33] <= 0;
			buffer[ 34] <= 0;
			buffer[ 35] <= 0;
			buffer[ 36] <= 0;
			buffer[ 37] <= 0;
			buffer[ 38] <= 0;
			buffer[ 39] <= 0;
			buffer[ 40] <= 0;
			buffer[ 41] <= 0;
			buffer[ 42] <= 0;
			buffer[ 43] <= 0;
			buffer[ 44] <= 0;
			buffer[ 45] <= 0;
			buffer[ 46] <= 0;
			buffer[ 47] <= 0;
			buffer[ 48] <= 0;
			buffer[ 49] <= 0;
			buffer[ 50] <= 0;
			buffer[ 51] <= 0;
			buffer[ 52] <= 0;
			buffer[ 53] <= 0;
			buffer[ 54] <= 0;
			buffer[ 55] <= 0;
			buffer[ 56] <= 0;
			buffer[ 57] <= 0;
			buffer[ 58] <= 0;
			buffer[ 59] <= 0;
			buffer[ 60] <= 0;
			buffer[ 61] <= 0;
			buffer[ 62] <= 0;
			buffer[ 63] <= 0;
			buffer[ 64] <= 0;
			buffer[ 65] <= 0;
			buffer[ 66] <= 0;
			buffer[ 67] <= 0;
			buffer[ 68] <= 0;
			buffer[ 69] <= 0;
			buffer[ 70] <= 0;
			buffer[ 71] <= 0;
			buffer[ 72] <= 0;
			buffer[ 73] <= 0;
			buffer[ 74] <= 0;
			buffer[ 75] <= 0;
			buffer[ 76] <= 0;
			buffer[ 77] <= 0;
			buffer[ 78] <= 0;
			buffer[ 79] <= 0;
			buffer[ 80] <= 0;
			buffer[ 81] <= 0;
			buffer[ 82] <= 0;
			buffer[ 83] <= 0;
			buffer[ 84] <= 0;
			buffer[ 85] <= 0;
			buffer[ 86] <= 0;
			buffer[ 87] <= 0;
			buffer[ 88] <= 0;
			buffer[ 89] <= 0;
			buffer[ 90] <= 0;
			buffer[ 91] <= 0;
			buffer[ 92] <= 0;
			buffer[ 93] <= 0;
			buffer[ 94] <= 0;
			buffer[ 95] <= 0;
			buffer[ 96] <= 0;
			buffer[ 97] <= 0;
			buffer[ 98] <= 0;
			buffer[ 99] <= 0;
			buffer[100] <= 0;
			buffer[101] <= 0;
			buffer[102] <= 0;
			buffer[103] <= 0;
			buffer[104] <= 0;
			buffer[105] <= 0;
			buffer[106] <= 0;
			buffer[107] <= 0;
			buffer[108] <= 0;
			buffer[109] <= 0;
			buffer[110] <= 0;
			buffer[111] <= 0;
			buffer[112] <= 0;
			buffer[113] <= 0;
			buffer[114] <= 0;
			buffer[115] <= 0;
			buffer[116] <= 0;
			buffer[117] <= 0;
			buffer[118] <= 0;
			buffer[119] <= 0;
			buffer[120] <= 0;
			buffer[121] <= 0;
			buffer[122] <= 0;
			buffer[123] <= 0;
			buffer[124] <= 0;
			buffer[125] <= 0;
			buffer[126] <= 0;
			buffer[127] <= 0;
			buffer[128] <= 0;
			buffer[129] <= 0;
			buffer[130] <= 0;
			buffer[131] <= 0;
			buffer[132] <= 0;
			buffer[133] <= 0;
			buffer[134] <= 0;
			buffer[135] <= 0;
			buffer[136] <= 0;
			buffer[137] <= 0;
			buffer[138] <= 0;
			buffer[139] <= 0;
			buffer[140] <= 0;
			buffer[141] <= 0;
			buffer[142] <= 0;
			buffer[143] <= 0;
			buffer[144] <= 0;
			buffer[145] <= 0;
			buffer[146] <= 0;
			buffer[147] <= 0;
			buffer[148] <= 0;
			buffer[149] <= 0;
			buffer[150] <= 0;
			buffer[151] <= 0;
			buffer[152] <= 0;
			buffer[153] <= 0;
			buffer[154] <= 0;
			buffer[155] <= 0;
			buffer[156] <= 0;
			buffer[157] <= 0;
			buffer[158] <= 0;
			buffer[159] <= 0;
			buffer[160] <= 0;
			buffer[161] <= 0;
			buffer[162] <= 0;
			buffer[163] <= 0;
			buffer[164] <= 0;
			buffer[165] <= 0;
			buffer[166] <= 0;
			buffer[167] <= 0;
			buffer[168] <= 0;
			buffer[169] <= 0;
			buffer[170] <= 0;
			buffer[171] <= 0;
			buffer[172] <= 0;
			buffer[173] <= 0;
			buffer[174] <= 0;
			buffer[175] <= 0;
			buffer[176] <= 0;
			buffer[177] <= 0;
			buffer[178] <= 0;
			buffer[179] <= 0;
			buffer[180] <= 0;
			buffer[181] <= 0;
			buffer[182] <= 0;
			buffer[183] <= 0;
			buffer[184] <= 0;
			buffer[185] <= 0;
			buffer[186] <= 0;
			buffer[187] <= 0;
			buffer[188] <= 0;
			buffer[189] <= 0;
			buffer[190] <= 0;
			buffer[191] <= 0;
			buffer[192] <= 0;
			buffer[193] <= 0;
			buffer[194] <= 0;
			buffer[195] <= 0;
			buffer[196] <= 0;
			buffer[197] <= 0;
			buffer[198] <= 0;
			buffer[199] <= 0;
			buffer[200] <= 0;
			buffer[201] <= 0;
			buffer[202] <= 0;
			buffer[203] <= 0;
			buffer[204] <= 0;
			buffer[205] <= 0;
			buffer[206] <= 0;
			buffer[207] <= 0;
			buffer[208] <= 0;
			buffer[209] <= 0;
			buffer[210] <= 0;
			buffer[211] <= 0;
			buffer[212] <= 0;
			buffer[213] <= 0;
			buffer[214] <= 0;
			buffer[215] <= 0;
			buffer[216] <= 0;
			buffer[217] <= 0;
			buffer[218] <= 0;
			buffer[219] <= 0;
			buffer[220] <= 0;
			buffer[221] <= 0;
			buffer[222] <= 0;
			buffer[223] <= 0;
			buffer[224] <= 0;
			buffer[225] <= 0;
			buffer[226] <= 0;
			buffer[227] <= 0;
			buffer[228] <= 0;
			buffer[229] <= 0;
			buffer[230] <= 0;
			buffer[231] <= 0;
			buffer[232] <= 0;
			buffer[233] <= 0;
			buffer[234] <= 0;
			buffer[235] <= 0;
			buffer[236] <= 0;
			buffer[237] <= 0;
			buffer[238] <= 0;
			buffer[239] <= 0;
			buffer[240] <= 0;
			buffer[241] <= 0;
			buffer[242] <= 0;
			buffer[243] <= 0;
			buffer[244] <= 0;
			buffer[245] <= 0;
			buffer[246] <= 0;
			buffer[247] <= 0;
			buffer[248] <= 0;
			buffer[249] <= 0;
			buffer[250] <= 0;
			buffer[251] <= 0;
			buffer[252] <= 0;
			buffer[253] <= 0;
			buffer[254] <= 0;
			buffer[255] <= 0;
		end else begin
			if (i_result_in_en) begin
				buffer[  0] <= i_data0;
				buffer[  1] <= i_data1;
				buffer[  2] <= i_data2;
				buffer[  3] <= i_data3;
				buffer[  4] <= i_data4;
				buffer[  5] <= i_data5;
				buffer[  6] <= i_data6;
				buffer[  7] <= i_data7;
				buffer[  8] <= i_data8;
				buffer[  9] <= i_data9;
				buffer[ 10] <= i_data10;
				buffer[ 11] <= i_data11;
				buffer[ 12] <= i_data12;
				buffer[ 13] <= i_data13;
				buffer[ 14] <= i_data14;
				buffer[ 15] <= i_data15;
				buffer[ 16] <= i_data16;
				buffer[ 17] <= i_data17;
				buffer[ 18] <= i_data18;
				buffer[ 19] <= i_data19;
				buffer[ 20] <= i_data20;
				buffer[ 21] <= i_data21;
				buffer[ 22] <= i_data22;
				buffer[ 23] <= i_data23;
				buffer[ 24] <= i_data24;
				buffer[ 25] <= i_data25;
				buffer[ 26] <= i_data26;
				buffer[ 27] <= i_data27;
				buffer[ 28] <= i_data28;
				buffer[ 29] <= i_data29;
				buffer[ 30] <= i_data30;
				buffer[ 31] <= i_data31;
				buffer[ 32] <= i_data32;
				buffer[ 33] <= i_data33;
				buffer[ 34] <= i_data34;
				buffer[ 35] <= i_data35;
				buffer[ 36] <= i_data36;
				buffer[ 37] <= i_data37;
				buffer[ 38] <= i_data38;
				buffer[ 39] <= i_data39;
				buffer[ 40] <= i_data40;
				buffer[ 41] <= i_data41;
				buffer[ 42] <= i_data42;
				buffer[ 43] <= i_data43;
				buffer[ 44] <= i_data44;
				buffer[ 45] <= i_data45;
				buffer[ 46] <= i_data46;
				buffer[ 47] <= i_data47;
				buffer[ 48] <= i_data48;
				buffer[ 49] <= i_data49;
				buffer[ 50] <= i_data50;
				buffer[ 51] <= i_data51;
				buffer[ 52] <= i_data52;
				buffer[ 53] <= i_data53;
				buffer[ 54] <= i_data54;
				buffer[ 55] <= i_data55;
				buffer[ 56] <= i_data56;
				buffer[ 57] <= i_data57;
				buffer[ 58] <= i_data58;
				buffer[ 59] <= i_data59;
				buffer[ 60] <= i_data60;
				buffer[ 61] <= i_data61;
				buffer[ 62] <= i_data62;
				buffer[ 63] <= i_data63;
				buffer[ 64] <= i_data64;
				buffer[ 65] <= i_data65;
				buffer[ 66] <= i_data66;
				buffer[ 67] <= i_data67;
				buffer[ 68] <= i_data68;
				buffer[ 69] <= i_data69;
				buffer[ 70] <= i_data70;
				buffer[ 71] <= i_data71;
				buffer[ 72] <= i_data72;
				buffer[ 73] <= i_data73;
				buffer[ 74] <= i_data74;
				buffer[ 75] <= i_data75;
				buffer[ 76] <= i_data76;
				buffer[ 77] <= i_data77;
				buffer[ 78] <= i_data78;
				buffer[ 79] <= i_data79;
				buffer[ 80] <= i_data80;
				buffer[ 81] <= i_data81;
				buffer[ 82] <= i_data82;
				buffer[ 83] <= i_data83;
				buffer[ 84] <= i_data84;
				buffer[ 85] <= i_data85;
				buffer[ 86] <= i_data86;
				buffer[ 87] <= i_data87;
				buffer[ 88] <= i_data88;
				buffer[ 89] <= i_data89;
				buffer[ 90] <= i_data90;
				buffer[ 91] <= i_data91;
				buffer[ 92] <= i_data92;
				buffer[ 93] <= i_data93;
				buffer[ 94] <= i_data94;
				buffer[ 95] <= i_data95;
				buffer[ 96] <= i_data96;
				buffer[ 97] <= i_data97;
				buffer[ 98] <= i_data98;
				buffer[ 99] <= i_data99;
				buffer[100] <= i_data100;
				buffer[101] <= i_data101;
				buffer[102] <= i_data102;
				buffer[103] <= i_data103;
				buffer[104] <= i_data104;
				buffer[105] <= i_data105;
				buffer[106] <= i_data106;
				buffer[107] <= i_data107;
				buffer[108] <= i_data108;
				buffer[109] <= i_data109;
				buffer[110] <= i_data110;
				buffer[111] <= i_data111;
				buffer[112] <= i_data112;
				buffer[113] <= i_data113;
				buffer[114] <= i_data114;
				buffer[115] <= i_data115;
				buffer[116] <= i_data116;
				buffer[117] <= i_data117;
				buffer[118] <= i_data118;
				buffer[119] <= i_data119;
				buffer[120] <= i_data120;
				buffer[121] <= i_data121;
				buffer[122] <= i_data122;
				buffer[123] <= i_data123;
				buffer[124] <= i_data124;
				buffer[125] <= i_data125;
				buffer[126] <= i_data126;
				buffer[127] <= i_data127;
				buffer[128] <= i_data128;
				buffer[129] <= i_data129;
				buffer[130] <= i_data130;
				buffer[131] <= i_data131;
				buffer[132] <= i_data132;
				buffer[133] <= i_data133;
				buffer[134] <= i_data134;
				buffer[135] <= i_data135;
				buffer[136] <= i_data136;
				buffer[137] <= i_data137;
				buffer[138] <= i_data138;
				buffer[139] <= i_data139;
				buffer[140] <= i_data140;
				buffer[141] <= i_data141;
				buffer[142] <= i_data142;
				buffer[143] <= i_data143;
				buffer[144] <= i_data144;
				buffer[145] <= i_data145;
				buffer[146] <= i_data146;
				buffer[147] <= i_data147;
				buffer[148] <= i_data148;
				buffer[149] <= i_data149;
				buffer[150] <= i_data150;
				buffer[151] <= i_data151;
				buffer[152] <= i_data152;
				buffer[153] <= i_data153;
				buffer[154] <= i_data154;
				buffer[155] <= i_data155;
				buffer[156] <= i_data156;
				buffer[157] <= i_data157;
				buffer[158] <= i_data158;
				buffer[159] <= i_data159;
				buffer[160] <= i_data160;
				buffer[161] <= i_data161;
				buffer[162] <= i_data162;
				buffer[163] <= i_data163;
				buffer[164] <= i_data164;
				buffer[165] <= i_data165;
				buffer[166] <= i_data166;
				buffer[167] <= i_data167;
				buffer[168] <= i_data168;
				buffer[169] <= i_data169;
				buffer[170] <= i_data170;
				buffer[171] <= i_data171;
				buffer[172] <= i_data172;
				buffer[173] <= i_data173;
				buffer[174] <= i_data174;
				buffer[175] <= i_data175;
				buffer[176] <= i_data176;
				buffer[177] <= i_data177;
				buffer[178] <= i_data178;
				buffer[179] <= i_data179;
				buffer[180] <= i_data180;
				buffer[181] <= i_data181;
				buffer[182] <= i_data182;
				buffer[183] <= i_data183;
				buffer[184] <= i_data184;
				buffer[185] <= i_data185;
				buffer[186] <= i_data186;
				buffer[187] <= i_data187;
				buffer[188] <= i_data188;
				buffer[189] <= i_data189;
				buffer[190] <= i_data190;
				buffer[191] <= i_data191;
				buffer[192] <= i_data192;
				buffer[193] <= i_data193;
				buffer[194] <= i_data194;
				buffer[195] <= i_data195;
				buffer[196] <= i_data196;
				buffer[197] <= i_data197;
				buffer[198] <= i_data198;
				buffer[199] <= i_data199;
				buffer[200] <= i_data200;
				buffer[201] <= i_data201;
				buffer[202] <= i_data202;
				buffer[203] <= i_data203;
				buffer[204] <= i_data204;
				buffer[205] <= i_data205;
				buffer[206] <= i_data206;
				buffer[207] <= i_data207;
				buffer[208] <= i_data208;
				buffer[209] <= i_data209;
				buffer[210] <= i_data210;
				buffer[211] <= i_data211;
				buffer[212] <= i_data212;
				buffer[213] <= i_data213;
				buffer[214] <= i_data214;
				buffer[215] <= i_data215;
				buffer[216] <= i_data216;
				buffer[217] <= i_data217;
				buffer[218] <= i_data218;
				buffer[219] <= i_data219;
				buffer[220] <= i_data220;
				buffer[221] <= i_data221;
				buffer[222] <= i_data222;
				buffer[223] <= i_data223;
				buffer[224] <= i_data224;
				buffer[225] <= i_data225;
				buffer[226] <= i_data226;
				buffer[227] <= i_data227;
				buffer[228] <= i_data228;
				buffer[229] <= i_data229;
				buffer[230] <= i_data230;
				buffer[231] <= i_data231;
				buffer[232] <= i_data232;
				buffer[233] <= i_data233;
				buffer[234] <= i_data234;
				buffer[235] <= i_data235;
				buffer[236] <= i_data236;
				buffer[237] <= i_data237;
				buffer[238] <= i_data238;
				buffer[239] <= i_data239;
				buffer[240] <= i_data240;
				buffer[241] <= i_data241;
				buffer[242] <= i_data242;
				buffer[243] <= i_data243;
				buffer[244] <= i_data244;
				buffer[245] <= i_data245;
				buffer[246] <= i_data246;
				buffer[247] <= i_data247;
				buffer[248] <= i_data248;
				buffer[249] <= i_data249;
				buffer[250] <= i_data250;
				buffer[251] <= i_data251;
				buffer[252] <= i_data252;
				buffer[253] <= i_data253;
				buffer[254] <= i_data254;
				buffer[255] <= i_data255;
			end
		end
	end

	assign o_data = i_result_out_en ? buffer[i_counter] : 0;


endmodule

// module result_buffer (
// 	input CLK,
// 	input !RSTN,
// 	input i_result_buffer_busy,
// 	input i_result_in_en,
// 	input i_result_out_en,
// 	input [7:0] i_counter,
// 	input [8191:0] i_data,
// 	output reg [31:0] o_data
// );

// 	reg [31:0] buffer [0:255];

// 	always @(posedge CLK) begin
// 		if (!RSTN) begin
// 			buffer[  0] <= 0;
// 			buffer[  1] <= 0;
// 			buffer[  2] <= 0;
// 			buffer[  3] <= 0;
// 			buffer[  4] <= 0;
// 			buffer[  5] <= 0;
// 			buffer[  6] <= 0;
// 			buffer[  7] <= 0;
// 			buffer[  8] <= 0;
// 			buffer[  9] <= 0;
// 			buffer[ 10] <= 0;
// 			buffer[ 11] <= 0;
// 			buffer[ 12] <= 0;
// 			buffer[ 13] <= 0;
// 			buffer[ 14] <= 0;
// 			buffer[ 15] <= 0;
// 			buffer[ 16] <= 0;
// 			buffer[ 17] <= 0;
// 			buffer[ 18] <= 0;
// 			buffer[ 19] <= 0;
// 			buffer[ 20] <= 0;
// 			buffer[ 21] <= 0;
// 			buffer[ 22] <= 0;
// 			buffer[ 23] <= 0;
// 			buffer[ 24] <= 0;
// 			buffer[ 25] <= 0;
// 			buffer[ 26] <= 0;
// 			buffer[ 27] <= 0;
// 			buffer[ 28] <= 0;
// 			buffer[ 29] <= 0;
// 			buffer[ 30] <= 0;
// 			buffer[ 31] <= 0;
// 			buffer[ 32] <= 0;
// 			buffer[ 33] <= 0;
// 			buffer[ 34] <= 0;
// 			buffer[ 35] <= 0;
// 			buffer[ 36] <= 0;
// 			buffer[ 37] <= 0;
// 			buffer[ 38] <= 0;
// 			buffer[ 39] <= 0;
// 			buffer[ 40] <= 0;
// 			buffer[ 41] <= 0;
// 			buffer[ 42] <= 0;
// 			buffer[ 43] <= 0;
// 			buffer[ 44] <= 0;
// 			buffer[ 45] <= 0;
// 			buffer[ 46] <= 0;
// 			buffer[ 47] <= 0;
// 			buffer[ 48] <= 0;
// 			buffer[ 49] <= 0;
// 			buffer[ 50] <= 0;
// 			buffer[ 51] <= 0;
// 			buffer[ 52] <= 0;
// 			buffer[ 53] <= 0;
// 			buffer[ 54] <= 0;
// 			buffer[ 55] <= 0;
// 			buffer[ 56] <= 0;
// 			buffer[ 57] <= 0;
// 			buffer[ 58] <= 0;
// 			buffer[ 59] <= 0;
// 			buffer[ 60] <= 0;
// 			buffer[ 61] <= 0;
// 			buffer[ 62] <= 0;
// 			buffer[ 63] <= 0;
// 			buffer[ 64] <= 0;
// 			buffer[ 65] <= 0;
// 			buffer[ 66] <= 0;
// 			buffer[ 67] <= 0;
// 			buffer[ 68] <= 0;
// 			buffer[ 69] <= 0;
// 			buffer[ 70] <= 0;
// 			buffer[ 71] <= 0;
// 			buffer[ 72] <= 0;
// 			buffer[ 73] <= 0;
// 			buffer[ 74] <= 0;
// 			buffer[ 75] <= 0;
// 			buffer[ 76] <= 0;
// 			buffer[ 77] <= 0;
// 			buffer[ 78] <= 0;
// 			buffer[ 79] <= 0;
// 			buffer[ 80] <= 0;
// 			buffer[ 81] <= 0;
// 			buffer[ 82] <= 0;
// 			buffer[ 83] <= 0;
// 			buffer[ 84] <= 0;
// 			buffer[ 85] <= 0;
// 			buffer[ 86] <= 0;
// 			buffer[ 87] <= 0;
// 			buffer[ 88] <= 0;
// 			buffer[ 89] <= 0;
// 			buffer[ 90] <= 0;
// 			buffer[ 91] <= 0;
// 			buffer[ 92] <= 0;
// 			buffer[ 93] <= 0;
// 			buffer[ 94] <= 0;
// 			buffer[ 95] <= 0;
// 			buffer[ 96] <= 0;
// 			buffer[ 97] <= 0;
// 			buffer[ 98] <= 0;
// 			buffer[ 99] <= 0;
// 			buffer[100] <= 0;
// 			buffer[101] <= 0;
// 			buffer[102] <= 0;
// 			buffer[103] <= 0;
// 			buffer[104] <= 0;
// 			buffer[105] <= 0;
// 			buffer[106] <= 0;
// 			buffer[107] <= 0;
// 			buffer[108] <= 0;
// 			buffer[109] <= 0;
// 			buffer[110] <= 0;
// 			buffer[111] <= 0;
// 			buffer[112] <= 0;
// 			buffer[113] <= 0;
// 			buffer[114] <= 0;
// 			buffer[115] <= 0;
// 			buffer[116] <= 0;
// 			buffer[117] <= 0;
// 			buffer[118] <= 0;
// 			buffer[119] <= 0;
// 			buffer[120] <= 0;
// 			buffer[121] <= 0;
// 			buffer[122] <= 0;
// 			buffer[123] <= 0;
// 			buffer[124] <= 0;
// 			buffer[125] <= 0;
// 			buffer[126] <= 0;
// 			buffer[127] <= 0;
// 			buffer[128] <= 0;
// 			buffer[129] <= 0;
// 			buffer[130] <= 0;
// 			buffer[131] <= 0;
// 			buffer[132] <= 0;
// 			buffer[133] <= 0;
// 			buffer[134] <= 0;
// 			buffer[135] <= 0;
// 			buffer[136] <= 0;
// 			buffer[137] <= 0;
// 			buffer[138] <= 0;
// 			buffer[139] <= 0;
// 			buffer[140] <= 0;
// 			buffer[141] <= 0;
// 			buffer[142] <= 0;
// 			buffer[143] <= 0;
// 			buffer[144] <= 0;
// 			buffer[145] <= 0;
// 			buffer[146] <= 0;
// 			buffer[147] <= 0;
// 			buffer[148] <= 0;
// 			buffer[149] <= 0;
// 			buffer[150] <= 0;
// 			buffer[151] <= 0;
// 			buffer[152] <= 0;
// 			buffer[153] <= 0;
// 			buffer[154] <= 0;
// 			buffer[155] <= 0;
// 			buffer[156] <= 0;
// 			buffer[157] <= 0;
// 			buffer[158] <= 0;
// 			buffer[159] <= 0;
// 			buffer[160] <= 0;
// 			buffer[161] <= 0;
// 			buffer[162] <= 0;
// 			buffer[163] <= 0;
// 			buffer[164] <= 0;
// 			buffer[165] <= 0;
// 			buffer[166] <= 0;
// 			buffer[167] <= 0;
// 			buffer[168] <= 0;
// 			buffer[169] <= 0;
// 			buffer[170] <= 0;
// 			buffer[171] <= 0;
// 			buffer[172] <= 0;
// 			buffer[173] <= 0;
// 			buffer[174] <= 0;
// 			buffer[175] <= 0;
// 			buffer[176] <= 0;
// 			buffer[177] <= 0;
// 			buffer[178] <= 0;
// 			buffer[179] <= 0;
// 			buffer[180] <= 0;
// 			buffer[181] <= 0;
// 			buffer[182] <= 0;
// 			buffer[183] <= 0;
// 			buffer[184] <= 0;
// 			buffer[185] <= 0;
// 			buffer[186] <= 0;
// 			buffer[187] <= 0;
// 			buffer[188] <= 0;
// 			buffer[189] <= 0;
// 			buffer[190] <= 0;
// 			buffer[191] <= 0;
// 			buffer[192] <= 0;
// 			buffer[193] <= 0;
// 			buffer[194] <= 0;
// 			buffer[195] <= 0;
// 			buffer[196] <= 0;
// 			buffer[197] <= 0;
// 			buffer[198] <= 0;
// 			buffer[199] <= 0;
// 			buffer[200] <= 0;
// 			buffer[201] <= 0;
// 			buffer[202] <= 0;
// 			buffer[203] <= 0;
// 			buffer[204] <= 0;
// 			buffer[205] <= 0;
// 			buffer[206] <= 0;
// 			buffer[207] <= 0;
// 			buffer[208] <= 0;
// 			buffer[209] <= 0;
// 			buffer[210] <= 0;
// 			buffer[211] <= 0;
// 			buffer[212] <= 0;
// 			buffer[213] <= 0;
// 			buffer[214] <= 0;
// 			buffer[215] <= 0;
// 			buffer[216] <= 0;
// 			buffer[217] <= 0;
// 			buffer[218] <= 0;
// 			buffer[219] <= 0;
// 			buffer[220] <= 0;
// 			buffer[221] <= 0;
// 			buffer[222] <= 0;
// 			buffer[223] <= 0;
// 			buffer[224] <= 0;
// 			buffer[225] <= 0;
// 			buffer[226] <= 0;
// 			buffer[227] <= 0;
// 			buffer[228] <= 0;
// 			buffer[229] <= 0;
// 			buffer[230] <= 0;
// 			buffer[231] <= 0;
// 			buffer[232] <= 0;
// 			buffer[233] <= 0;
// 			buffer[234] <= 0;
// 			buffer[235] <= 0;
// 			buffer[236] <= 0;
// 			buffer[237] <= 0;
// 			buffer[238] <= 0;
// 			buffer[239] <= 0;
// 			buffer[240] <= 0;
// 			buffer[241] <= 0;
// 			buffer[242] <= 0;
// 			buffer[243] <= 0;
// 			buffer[244] <= 0;
// 			buffer[245] <= 0;
// 			buffer[246] <= 0;
// 			buffer[247] <= 0;
// 			buffer[248] <= 0;
// 			buffer[249] <= 0;
// 			buffer[250] <= 0;
// 			buffer[251] <= 0;
// 			buffer[252] <= 0;
// 			buffer[253] <= 0;
// 			buffer[254] <= 0;
// 			buffer[255] <= 0;
// 		end else begin
// 			if (i_result_buffer_busy) begin
// 				if (i_result_in_en) begin
// 				buffer[  0] <= i_data[8191:8160];
// 				buffer[  1] <= i_data[8159:8128];
// 				buffer[  2] <= i_data[8127:8096];
// 				buffer[  3] <= i_data[8095:8064];
// 				buffer[  4] <= i_data[8063:8032];
// 				buffer[  5] <= i_data[8031:8000];
// 				buffer[  6] <= i_data[7999:7968];
// 				buffer[  7] <= i_data[7967:7936];
// 				buffer[  8] <= i_data[7935:7904];
// 				buffer[  9] <= i_data[7903:7872];
// 				buffer[ 10] <= i_data[7871:7840];
// 				buffer[ 11] <= i_data[7839:7808];
// 				buffer[ 12] <= i_data[7807:7776];
// 				buffer[ 13] <= i_data[7775:7744];
// 				buffer[ 14] <= i_data[7743:7712];
// 				buffer[ 15] <= i_data[7711:7680];
// 				buffer[ 16] <= i_data[7679:7648];
// 				buffer[ 17] <= i_data[7647:7616];
// 				buffer[ 18] <= i_data[7615:7584];
// 				buffer[ 19] <= i_data[7583:7552];
// 				buffer[ 20] <= i_data[7551:7520];
// 				buffer[ 21] <= i_data[7519:7488];
// 				buffer[ 22] <= i_data[7487:7456];
// 				buffer[ 23] <= i_data[7455:7424];
// 				buffer[ 24] <= i_data[7423:7392];
// 				buffer[ 25] <= i_data[7391:7360];
// 				buffer[ 26] <= i_data[7359:7328];
// 				buffer[ 27] <= i_data[7327:7296];
// 				buffer[ 28] <= i_data[7295:7264];
// 				buffer[ 29] <= i_data[7263:7232];
// 				buffer[ 30] <= i_data[7231:7200];
// 				buffer[ 31] <= i_data[7199:7168];
// 				buffer[ 32] <= i_data[7167:7136];
// 				buffer[ 33] <= i_data[7135:7104];
// 				buffer[ 34] <= i_data[7103:7072];
// 				buffer[ 35] <= i_data[7071:7040];
// 				buffer[ 36] <= i_data[7039:7008];
// 				buffer[ 37] <= i_data[7007:6976];
// 				buffer[ 38] <= i_data[6975:6944];
// 				buffer[ 39] <= i_data[6943:6912];
// 				buffer[ 40] <= i_data[6911:6880];
// 				buffer[ 41] <= i_data[6879:6848];
// 				buffer[ 42] <= i_data[6847:6816];
// 				buffer[ 43] <= i_data[6815:6784];
// 				buffer[ 44] <= i_data[6783:6752];
// 				buffer[ 45] <= i_data[6751:6720];
// 				buffer[ 46] <= i_data[6719:6688];
// 				buffer[ 47] <= i_data[6687:6656];
// 				buffer[ 48] <= i_data[6655:6624];
// 				buffer[ 49] <= i_data[6623:6592];
// 				buffer[ 50] <= i_data[6591:6560];
// 				buffer[ 51] <= i_data[6559:6528];
// 				buffer[ 52] <= i_data[6527:6496];
// 				buffer[ 53] <= i_data[6495:6464];
// 				buffer[ 54] <= i_data[6463:6432];
// 				buffer[ 55] <= i_data[6431:6400];
// 				buffer[ 56] <= i_data[6399:6368];
// 				buffer[ 57] <= i_data[6367:6336];
// 				buffer[ 58] <= i_data[6335:6304];
// 				buffer[ 59] <= i_data[6303:6272];
// 				buffer[ 60] <= i_data[6271:6240];
// 				buffer[ 61] <= i_data[6239:6208];
// 				buffer[ 62] <= i_data[6207:6176];
// 				buffer[ 63] <= i_data[6175:6144];
// 				buffer[ 64] <= i_data[6143:6112];
// 				buffer[ 65] <= i_data[6111:6080];
// 				buffer[ 66] <= i_data[6079:6048];
// 				buffer[ 67] <= i_data[6047:6016];
// 				buffer[ 68] <= i_data[6015:5984];
// 				buffer[ 69] <= i_data[5983:5952];
// 				buffer[ 70] <= i_data[5951:5920];
// 				buffer[ 71] <= i_data[5919:5888];
// 				buffer[ 72] <= i_data[5887:5856];
// 				buffer[ 73] <= i_data[5855:5824];
// 				buffer[ 74] <= i_data[5823:5792];
// 				buffer[ 75] <= i_data[5791:5760];
// 				buffer[ 76] <= i_data[5759:5728];
// 				buffer[ 77] <= i_data[5727:5696];
// 				buffer[ 78] <= i_data[5695:5664];
// 				buffer[ 79] <= i_data[5663:5632];
// 				buffer[ 80] <= i_data[5631:5600];
// 				buffer[ 81] <= i_data[5599:5568];
// 				buffer[ 82] <= i_data[5567:5536];
// 				buffer[ 83] <= i_data[5535:5504];
// 				buffer[ 84] <= i_data[5503:5472];
// 				buffer[ 85] <= i_data[5471:5440];
// 				buffer[ 86] <= i_data[5439:5408];
// 				buffer[ 87] <= i_data[5407:5376];
// 				buffer[ 88] <= i_data[5375:5344];
// 				buffer[ 89] <= i_data[5343:5312];
// 				buffer[ 90] <= i_data[5311:5280];
// 				buffer[ 91] <= i_data[5279:5248];
// 				buffer[ 92] <= i_data[5247:5216];
// 				buffer[ 93] <= i_data[5215:5184];
// 				buffer[ 94] <= i_data[5183:5152];
// 				buffer[ 95] <= i_data[5151:5120];
// 				buffer[ 96] <= i_data[5119:5088];
// 				buffer[ 97] <= i_data[5087:5056];
// 				buffer[ 98] <= i_data[5055:5024];
// 				buffer[ 99] <= i_data[5023:4992];
// 				buffer[100] <= i_data[4991:4960];
// 				buffer[101] <= i_data[4959:4928];
// 				buffer[102] <= i_data[4927:4896];
// 				buffer[103] <= i_data[4895:4864];
// 				buffer[104] <= i_data[4863:4832];
// 				buffer[105] <= i_data[4831:4800];
// 				buffer[106] <= i_data[4799:4768];
// 				buffer[107] <= i_data[4767:4736];
// 				buffer[108] <= i_data[4735:4704];
// 				buffer[109] <= i_data[4703:4672];
// 				buffer[110] <= i_data[4671:4640];
// 				buffer[111] <= i_data[4639:4608];
// 				buffer[112] <= i_data[4607:4576];
// 				buffer[113] <= i_data[4575:4544];
// 				buffer[114] <= i_data[4543:4512];
// 				buffer[115] <= i_data[4511:4480];
// 				buffer[116] <= i_data[4479:4448];
// 				buffer[117] <= i_data[4447:4416];
// 				buffer[118] <= i_data[4415:4384];
// 				buffer[119] <= i_data[4383:4352];
// 				buffer[120] <= i_data[4351:4320];
// 				buffer[121] <= i_data[4319:4288];
// 				buffer[122] <= i_data[4287:4256];
// 				buffer[123] <= i_data[4255:4224];
// 				buffer[124] <= i_data[4223:4192];
// 				buffer[125] <= i_data[4191:4160];
// 				buffer[126] <= i_data[4159:4128];
// 				buffer[127] <= i_data[4127:4096];
// 				buffer[128] <= i_data[4095:4064];
// 				buffer[129] <= i_data[4063:4032];
// 				buffer[130] <= i_data[4031:4000];
// 				buffer[131] <= i_data[3999:3968];
// 				buffer[132] <= i_data[3967:3936];
// 				buffer[133] <= i_data[3935:3904];
// 				buffer[134] <= i_data[3903:3872];
// 				buffer[135] <= i_data[3871:3840];
// 				buffer[136] <= i_data[3839:3808];
// 				buffer[137] <= i_data[3807:3776];
// 				buffer[138] <= i_data[3775:3744];
// 				buffer[139] <= i_data[3743:3712];
// 				buffer[140] <= i_data[3711:3680];
// 				buffer[141] <= i_data[3679:3648];
// 				buffer[142] <= i_data[3647:3616];
// 				buffer[143] <= i_data[3615:3584];
// 				buffer[144] <= i_data[3583:3552];
// 				buffer[145] <= i_data[3551:3520];
// 				buffer[146] <= i_data[3519:3488];
// 				buffer[147] <= i_data[3487:3456];
// 				buffer[148] <= i_data[3455:3424];
// 				buffer[149] <= i_data[3423:3392];
// 				buffer[150] <= i_data[3391:3360];
// 				buffer[151] <= i_data[3359:3328];
// 				buffer[152] <= i_data[3327:3296];
// 				buffer[153] <= i_data[3295:3264];
// 				buffer[154] <= i_data[3263:3232];
// 				buffer[155] <= i_data[3231:3200];
// 				buffer[156] <= i_data[3199:3168];
// 				buffer[157] <= i_data[3167:3136];
// 				buffer[158] <= i_data[3135:3104];
// 				buffer[159] <= i_data[3103:3072];
// 				buffer[160] <= i_data[3071:3040];
// 				buffer[161] <= i_data[3039:3008];
// 				buffer[162] <= i_data[3007:2976];
// 				buffer[163] <= i_data[2975:2944];
// 				buffer[164] <= i_data[2943:2912];
// 				buffer[165] <= i_data[2911:2880];
// 				buffer[166] <= i_data[2879:2848];
// 				buffer[167] <= i_data[2847:2816];
// 				buffer[168] <= i_data[2815:2784];
// 				buffer[169] <= i_data[2783:2752];
// 				buffer[170] <= i_data[2751:2720];
// 				buffer[171] <= i_data[2719:2688];
// 				buffer[172] <= i_data[2687:2656];
// 				buffer[173] <= i_data[2655:2624];
// 				buffer[174] <= i_data[2623:2592];
// 				buffer[175] <= i_data[2591:2560];
// 				buffer[176] <= i_data[2559:2528];
// 				buffer[177] <= i_data[2527:2496];
// 				buffer[178] <= i_data[2495:2464];
// 				buffer[179] <= i_data[2463:2432];
// 				buffer[180] <= i_data[2431:2400];
// 				buffer[181] <= i_data[2399:2368];
// 				buffer[182] <= i_data[2367:2336];
// 				buffer[183] <= i_data[2335:2304];
// 				buffer[184] <= i_data[2303:2272];
// 				buffer[185] <= i_data[2271:2240];
// 				buffer[186] <= i_data[2239:2208];
// 				buffer[187] <= i_data[2207:2176];
// 				buffer[188] <= i_data[2175:2144];
// 				buffer[189] <= i_data[2143:2112];
// 				buffer[190] <= i_data[2111:2080];
// 				buffer[191] <= i_data[2079:2048];
// 				buffer[192] <= i_data[2047:2016];
// 				buffer[193] <= i_data[2015:1984];
// 				buffer[194] <= i_data[1983:1952];
// 				buffer[195] <= i_data[1951:1920];
// 				buffer[196] <= i_data[1919:1888];
// 				buffer[197] <= i_data[1887:1856];
// 				buffer[198] <= i_data[1855:1824];
// 				buffer[199] <= i_data[1823:1792];
// 				buffer[200] <= i_data[1791:1760];
// 				buffer[201] <= i_data[1759:1728];
// 				buffer[202] <= i_data[1727:1696];
// 				buffer[203] <= i_data[1695:1664];
// 				buffer[204] <= i_data[1663:1632];
// 				buffer[205] <= i_data[1631:1600];
// 				buffer[206] <= i_data[1599:1568];
// 				buffer[207] <= i_data[1567:1536];
// 				buffer[208] <= i_data[1535:1504];
// 				buffer[209] <= i_data[1503:1472];
// 				buffer[210] <= i_data[1471:1440];
// 				buffer[211] <= i_data[1439:1408];
// 				buffer[212] <= i_data[1407:1376];
// 				buffer[213] <= i_data[1375:1344];
// 				buffer[214] <= i_data[1343:1312];
// 				buffer[215] <= i_data[1311:1280];
// 				buffer[216] <= i_data[1279:1248];
// 				buffer[217] <= i_data[1247:1216];
// 				buffer[218] <= i_data[1215:1184];
// 				buffer[219] <= i_data[1183:1152];
// 				buffer[220] <= i_data[1151:1120];
// 				buffer[221] <= i_data[1119:1088];
// 				buffer[222] <= i_data[1087:1056];
// 				buffer[223] <= i_data[1055:1024];
// 				buffer[224] <= i_data[1023:992];
// 				buffer[225] <= i_data[991:960];
// 				buffer[226] <= i_data[959:928];
// 				buffer[227] <= i_data[927:896];
// 				buffer[228] <= i_data[895:864];
// 				buffer[229] <= i_data[863:832];
// 				buffer[230] <= i_data[831:800];
// 				buffer[231] <= i_data[799:768];
// 				buffer[232] <= i_data[767:736];
// 				buffer[233] <= i_data[735:704];
// 				buffer[234] <= i_data[703:672];
// 				buffer[235] <= i_data[671:640];
// 				buffer[236] <= i_data[639:608];
// 				buffer[237] <= i_data[607:576];
// 				buffer[238] <= i_data[575:544];
// 				buffer[239] <= i_data[543:512];
// 				buffer[240] <= i_data[511:480];
// 				buffer[241] <= i_data[479:448];
// 				buffer[242] <= i_data[447:416];
// 				buffer[243] <= i_data[415:384];
// 				buffer[244] <= i_data[383:352];
// 				buffer[245] <= i_data[351:320];
// 				buffer[246] <= i_data[319:288];
// 				buffer[247] <= i_data[287:256];
// 				buffer[248] <= i_data[255:224];
// 				buffer[249] <= i_data[223:192];
// 				buffer[250] <= i_data[191:160];
// 				buffer[251] <= i_data[159:128];
// 				buffer[252] <= i_data[127:96];
// 				buffer[253] <= i_data[95:64];
// 				buffer[254] <= i_data[63:32];
// 				buffer[255] <= i_data[31:0];
// 				end
// 			end else begin 
// 				buffer[  0] <= 0;
// 				buffer[  1] <= 0;
// 				buffer[  2] <= 0;
// 				buffer[  3] <= 0;
// 				buffer[  4] <= 0;
// 				buffer[  5] <= 0;
// 				buffer[  6] <= 0;
// 				buffer[  7] <= 0;
// 				buffer[  8] <= 0;
// 				buffer[  9] <= 0;
// 				buffer[ 10] <= 0;
// 				buffer[ 11] <= 0;
// 				buffer[ 12] <= 0;
// 				buffer[ 13] <= 0;
// 				buffer[ 14] <= 0;
// 				buffer[ 15] <= 0;
// 				buffer[ 16] <= 0;
// 				buffer[ 17] <= 0;
// 				buffer[ 18] <= 0;
// 				buffer[ 19] <= 0;
// 				buffer[ 20] <= 0;
// 				buffer[ 21] <= 0;
// 				buffer[ 22] <= 0;
// 				buffer[ 23] <= 0;
// 				buffer[ 24] <= 0;
// 				buffer[ 25] <= 0;
// 				buffer[ 26] <= 0;
// 				buffer[ 27] <= 0;
// 				buffer[ 28] <= 0;
// 				buffer[ 29] <= 0;
// 				buffer[ 30] <= 0;
// 				buffer[ 31] <= 0;
// 				buffer[ 32] <= 0;
// 				buffer[ 33] <= 0;
// 				buffer[ 34] <= 0;
// 				buffer[ 35] <= 0;
// 				buffer[ 36] <= 0;
// 				buffer[ 37] <= 0;
// 				buffer[ 38] <= 0;
// 				buffer[ 39] <= 0;
// 				buffer[ 40] <= 0;
// 				buffer[ 41] <= 0;
// 				buffer[ 42] <= 0;
// 				buffer[ 43] <= 0;
// 				buffer[ 44] <= 0;
// 				buffer[ 45] <= 0;
// 				buffer[ 46] <= 0;
// 				buffer[ 47] <= 0;
// 				buffer[ 48] <= 0;
// 				buffer[ 49] <= 0;
// 				buffer[ 50] <= 0;
// 				buffer[ 51] <= 0;
// 				buffer[ 52] <= 0;
// 				buffer[ 53] <= 0;
// 				buffer[ 54] <= 0;
// 				buffer[ 55] <= 0;
// 				buffer[ 56] <= 0;
// 				buffer[ 57] <= 0;
// 				buffer[ 58] <= 0;
// 				buffer[ 59] <= 0;
// 				buffer[ 60] <= 0;
// 				buffer[ 61] <= 0;
// 				buffer[ 62] <= 0;
// 				buffer[ 63] <= 0;
// 				buffer[ 64] <= 0;
// 				buffer[ 65] <= 0;
// 				buffer[ 66] <= 0;
// 				buffer[ 67] <= 0;
// 				buffer[ 68] <= 0;
// 				buffer[ 69] <= 0;
// 				buffer[ 70] <= 0;
// 				buffer[ 71] <= 0;
// 				buffer[ 72] <= 0;
// 				buffer[ 73] <= 0;
// 				buffer[ 74] <= 0;
// 				buffer[ 75] <= 0;
// 				buffer[ 76] <= 0;
// 				buffer[ 77] <= 0;
// 				buffer[ 78] <= 0;
// 				buffer[ 79] <= 0;
// 				buffer[ 80] <= 0;
// 				buffer[ 81] <= 0;
// 				buffer[ 82] <= 0;
// 				buffer[ 83] <= 0;
// 				buffer[ 84] <= 0;
// 				buffer[ 85] <= 0;
// 				buffer[ 86] <= 0;
// 				buffer[ 87] <= 0;
// 				buffer[ 88] <= 0;
// 				buffer[ 89] <= 0;
// 				buffer[ 90] <= 0;
// 				buffer[ 91] <= 0;
// 				buffer[ 92] <= 0;
// 				buffer[ 93] <= 0;
// 				buffer[ 94] <= 0;
// 				buffer[ 95] <= 0;
// 				buffer[ 96] <= 0;
// 				buffer[ 97] <= 0;
// 				buffer[ 98] <= 0;
// 				buffer[ 99] <= 0;
// 				buffer[100] <= 0;
// 				buffer[101] <= 0;
// 				buffer[102] <= 0;
// 				buffer[103] <= 0;
// 				buffer[104] <= 0;
// 				buffer[105] <= 0;
// 				buffer[106] <= 0;
// 				buffer[107] <= 0;
// 				buffer[108] <= 0;
// 				buffer[109] <= 0;
// 				buffer[110] <= 0;
// 				buffer[111] <= 0;
// 				buffer[112] <= 0;
// 				buffer[113] <= 0;
// 				buffer[114] <= 0;
// 				buffer[115] <= 0;
// 				buffer[116] <= 0;
// 				buffer[117] <= 0;
// 				buffer[118] <= 0;
// 				buffer[119] <= 0;
// 				buffer[120] <= 0;
// 				buffer[121] <= 0;
// 				buffer[122] <= 0;
// 				buffer[123] <= 0;
// 				buffer[124] <= 0;
// 				buffer[125] <= 0;
// 				buffer[126] <= 0;
// 				buffer[127] <= 0;
// 				buffer[128] <= 0;
// 				buffer[129] <= 0;
// 				buffer[130] <= 0;
// 				buffer[131] <= 0;
// 				buffer[132] <= 0;
// 				buffer[133] <= 0;
// 				buffer[134] <= 0;
// 				buffer[135] <= 0;
// 				buffer[136] <= 0;
// 				buffer[137] <= 0;
// 				buffer[138] <= 0;
// 				buffer[139] <= 0;
// 				buffer[140] <= 0;
// 				buffer[141] <= 0;
// 				buffer[142] <= 0;
// 				buffer[143] <= 0;
// 				buffer[144] <= 0;
// 				buffer[145] <= 0;
// 				buffer[146] <= 0;
// 				buffer[147] <= 0;
// 				buffer[148] <= 0;
// 				buffer[149] <= 0;
// 				buffer[150] <= 0;
// 				buffer[151] <= 0;
// 				buffer[152] <= 0;
// 				buffer[153] <= 0;
// 				buffer[154] <= 0;
// 				buffer[155] <= 0;
// 				buffer[156] <= 0;
// 				buffer[157] <= 0;
// 				buffer[158] <= 0;
// 				buffer[159] <= 0;
// 				buffer[160] <= 0;
// 				buffer[161] <= 0;
// 				buffer[162] <= 0;
// 				buffer[163] <= 0;
// 				buffer[164] <= 0;
// 				buffer[165] <= 0;
// 				buffer[166] <= 0;
// 				buffer[167] <= 0;
// 				buffer[168] <= 0;
// 				buffer[169] <= 0;
// 				buffer[170] <= 0;
// 				buffer[171] <= 0;
// 				buffer[172] <= 0;
// 				buffer[173] <= 0;
// 				buffer[174] <= 0;
// 				buffer[175] <= 0;
// 				buffer[176] <= 0;
// 				buffer[177] <= 0;
// 				buffer[178] <= 0;
// 				buffer[179] <= 0;
// 				buffer[180] <= 0;
// 				buffer[181] <= 0;
// 				buffer[182] <= 0;
// 				buffer[183] <= 0;
// 				buffer[184] <= 0;
// 				buffer[185] <= 0;
// 				buffer[186] <= 0;
// 				buffer[187] <= 0;
// 				buffer[188] <= 0;
// 				buffer[189] <= 0;
// 				buffer[190] <= 0;
// 				buffer[191] <= 0;
// 				buffer[192] <= 0;
// 				buffer[193] <= 0;
// 				buffer[194] <= 0;
// 				buffer[195] <= 0;
// 				buffer[196] <= 0;
// 				buffer[197] <= 0;
// 				buffer[198] <= 0;
// 				buffer[199] <= 0;
// 				buffer[200] <= 0;
// 				buffer[201] <= 0;
// 				buffer[202] <= 0;
// 				buffer[203] <= 0;
// 				buffer[204] <= 0;
// 				buffer[205] <= 0;
// 				buffer[206] <= 0;
// 				buffer[207] <= 0;
// 				buffer[208] <= 0;
// 				buffer[209] <= 0;
// 				buffer[210] <= 0;
// 				buffer[211] <= 0;
// 				buffer[212] <= 0;
// 				buffer[213] <= 0;
// 				buffer[214] <= 0;
// 				buffer[215] <= 0;
// 				buffer[216] <= 0;
// 				buffer[217] <= 0;
// 				buffer[218] <= 0;
// 				buffer[219] <= 0;
// 				buffer[220] <= 0;
// 				buffer[221] <= 0;
// 				buffer[222] <= 0;
// 				buffer[223] <= 0;
// 				buffer[224] <= 0;
// 				buffer[225] <= 0;
// 				buffer[226] <= 0;
// 				buffer[227] <= 0;
// 				buffer[228] <= 0;
// 				buffer[229] <= 0;
// 				buffer[230] <= 0;
// 				buffer[231] <= 0;
// 				buffer[232] <= 0;
// 				buffer[233] <= 0;
// 				buffer[234] <= 0;
// 				buffer[235] <= 0;
// 				buffer[236] <= 0;
// 				buffer[237] <= 0;
// 				buffer[238] <= 0;
// 				buffer[239] <= 0;
// 				buffer[240] <= 0;
// 				buffer[241] <= 0;
// 				buffer[242] <= 0;
// 				buffer[243] <= 0;
// 				buffer[244] <= 0;
// 				buffer[245] <= 0;
// 				buffer[246] <= 0;
// 				buffer[247] <= 0;
// 				buffer[248] <= 0;
// 				buffer[249] <= 0;
// 				buffer[250] <= 0;
// 				buffer[251] <= 0;
// 				buffer[252] <= 0;
// 				buffer[253] <= 0;
// 				buffer[254] <= 0;
// 				buffer[255] <= 0;
// 			end
// 		end
// 	end

// 	always @(*) begin
// 		if (!RSTN) begin
// 			o_data <= 0;
// 		end else begin
// 			if (i_result_out_en) begin
// 				o_data <= buffer[i_counter];
// 			end else begin
// 				o_data <= 0;
// 			end
// 		end
// 	end

// endmodule