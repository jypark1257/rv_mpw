module activation_buffer (
	input i_clk,
	input i_rst,
	input i_activation_in_en,
	input i_activation_out_en,
	input [7:0] i_counter,
	input [31:0] i_data,
	output reg [287:0] o_data
);

	reg [7:0] buffer [0:287];

	always @(posedge i_clk) begin
		if(i_rst) begin
			buffer[  0] <= 0;
			buffer[  1] <= 0;
			buffer[  2] <= 0;
			buffer[  3] <= 0;
			buffer[  4] <= 0;
			buffer[  5] <= 0;
			buffer[  6] <= 0;
			buffer[  7] <= 0;
			buffer[  8] <= 0;
			buffer[  9] <= 0;
			buffer[ 10] <= 0;
			buffer[ 11] <= 0;
			buffer[ 12] <= 0;
			buffer[ 13] <= 0;
			buffer[ 14] <= 0;
			buffer[ 15] <= 0;
			buffer[ 16] <= 0;
			buffer[ 17] <= 0;
			buffer[ 18] <= 0;
			buffer[ 19] <= 0;
			buffer[ 20] <= 0;
			buffer[ 21] <= 0;
			buffer[ 22] <= 0;
			buffer[ 23] <= 0;
			buffer[ 24] <= 0;
			buffer[ 25] <= 0;
			buffer[ 26] <= 0;
			buffer[ 27] <= 0;
			buffer[ 28] <= 0;
			buffer[ 29] <= 0;
			buffer[ 30] <= 0;
			buffer[ 31] <= 0;
			buffer[ 32] <= 0;
			buffer[ 33] <= 0;
			buffer[ 34] <= 0;
			buffer[ 35] <= 0;
			buffer[ 36] <= 0;
			buffer[ 37] <= 0;
			buffer[ 38] <= 0;
			buffer[ 39] <= 0;
			buffer[ 40] <= 0;
			buffer[ 41] <= 0;
			buffer[ 42] <= 0;
			buffer[ 43] <= 0;
			buffer[ 44] <= 0;
			buffer[ 45] <= 0;
			buffer[ 46] <= 0;
			buffer[ 47] <= 0;
			buffer[ 48] <= 0;
			buffer[ 49] <= 0;
			buffer[ 50] <= 0;
			buffer[ 51] <= 0;
			buffer[ 52] <= 0;
			buffer[ 53] <= 0;
			buffer[ 54] <= 0;
			buffer[ 55] <= 0;
			buffer[ 56] <= 0;
			buffer[ 57] <= 0;
			buffer[ 58] <= 0;
			buffer[ 59] <= 0;
			buffer[ 60] <= 0;
			buffer[ 61] <= 0;
			buffer[ 62] <= 0;
			buffer[ 63] <= 0;
			buffer[ 64] <= 0;
			buffer[ 65] <= 0;
			buffer[ 66] <= 0;
			buffer[ 67] <= 0;
			buffer[ 68] <= 0;
			buffer[ 69] <= 0;
			buffer[ 70] <= 0;
			buffer[ 71] <= 0;
			buffer[ 72] <= 0;
			buffer[ 73] <= 0;
			buffer[ 74] <= 0;
			buffer[ 75] <= 0;
			buffer[ 76] <= 0;
			buffer[ 77] <= 0;
			buffer[ 78] <= 0;
			buffer[ 79] <= 0;
			buffer[ 80] <= 0;
			buffer[ 81] <= 0;
			buffer[ 82] <= 0;
			buffer[ 83] <= 0;
			buffer[ 84] <= 0;
			buffer[ 85] <= 0;
			buffer[ 86] <= 0;
			buffer[ 87] <= 0;
			buffer[ 88] <= 0;
			buffer[ 89] <= 0;
			buffer[ 90] <= 0;
			buffer[ 91] <= 0;
			buffer[ 92] <= 0;
			buffer[ 93] <= 0;
			buffer[ 94] <= 0;
			buffer[ 95] <= 0;
			buffer[ 96] <= 0;
			buffer[ 97] <= 0;
			buffer[ 98] <= 0;
			buffer[ 99] <= 0;
			buffer[100] <= 0;
			buffer[101] <= 0;
			buffer[102] <= 0;
			buffer[103] <= 0;
			buffer[104] <= 0;
			buffer[105] <= 0;
			buffer[106] <= 0;
			buffer[107] <= 0;
			buffer[108] <= 0;
			buffer[109] <= 0;
			buffer[110] <= 0;
			buffer[111] <= 0;
			buffer[112] <= 0;
			buffer[113] <= 0;
			buffer[114] <= 0;
			buffer[115] <= 0;
			buffer[116] <= 0;
			buffer[117] <= 0;
			buffer[118] <= 0;
			buffer[119] <= 0;
			buffer[120] <= 0;
			buffer[121] <= 0;
			buffer[122] <= 0;
			buffer[123] <= 0;
			buffer[124] <= 0;
			buffer[125] <= 0;
			buffer[126] <= 0;
			buffer[127] <= 0;
			buffer[128] <= 0;
			buffer[129] <= 0;
			buffer[130] <= 0;
			buffer[131] <= 0;
			buffer[132] <= 0;
			buffer[133] <= 0;
			buffer[134] <= 0;
			buffer[135] <= 0;
			buffer[136] <= 0;
			buffer[137] <= 0;
			buffer[138] <= 0;
			buffer[139] <= 0;
			buffer[140] <= 0;
			buffer[141] <= 0;
			buffer[142] <= 0;
			buffer[143] <= 0;
			buffer[144] <= 0;
			buffer[145] <= 0;
			buffer[146] <= 0;
			buffer[147] <= 0;
			buffer[148] <= 0;
			buffer[149] <= 0;
			buffer[150] <= 0;
			buffer[151] <= 0;
			buffer[152] <= 0;
			buffer[153] <= 0;
			buffer[154] <= 0;
			buffer[155] <= 0;
			buffer[156] <= 0;
			buffer[157] <= 0;
			buffer[158] <= 0;
			buffer[159] <= 0;
			buffer[160] <= 0;
			buffer[161] <= 0;
			buffer[162] <= 0;
			buffer[163] <= 0;
			buffer[164] <= 0;
			buffer[165] <= 0;
			buffer[166] <= 0;
			buffer[167] <= 0;
			buffer[168] <= 0;
			buffer[169] <= 0;
			buffer[170] <= 0;
			buffer[171] <= 0;
			buffer[172] <= 0;
			buffer[173] <= 0;
			buffer[174] <= 0;
			buffer[175] <= 0;
			buffer[176] <= 0;
			buffer[177] <= 0;
			buffer[178] <= 0;
			buffer[179] <= 0;
			buffer[180] <= 0;
			buffer[181] <= 0;
			buffer[182] <= 0;
			buffer[183] <= 0;
			buffer[184] <= 0;
			buffer[185] <= 0;
			buffer[186] <= 0;
			buffer[187] <= 0;
			buffer[188] <= 0;
			buffer[189] <= 0;
			buffer[190] <= 0;
			buffer[191] <= 0;
			buffer[192] <= 0;
			buffer[193] <= 0;
			buffer[194] <= 0;
			buffer[195] <= 0;
			buffer[196] <= 0;
			buffer[197] <= 0;
			buffer[198] <= 0;
			buffer[199] <= 0;
			buffer[200] <= 0;
			buffer[201] <= 0;
			buffer[202] <= 0;
			buffer[203] <= 0;
			buffer[204] <= 0;
			buffer[205] <= 0;
			buffer[206] <= 0;
			buffer[207] <= 0;
			buffer[208] <= 0;
			buffer[209] <= 0;
			buffer[210] <= 0;
			buffer[211] <= 0;
			buffer[212] <= 0;
			buffer[213] <= 0;
			buffer[214] <= 0;
			buffer[215] <= 0;
			buffer[216] <= 0;
			buffer[217] <= 0;
			buffer[218] <= 0;
			buffer[219] <= 0;
			buffer[220] <= 0;
			buffer[221] <= 0;
			buffer[222] <= 0;
			buffer[223] <= 0;
			buffer[224] <= 0;
			buffer[225] <= 0;
			buffer[226] <= 0;
			buffer[227] <= 0;
			buffer[228] <= 0;
			buffer[229] <= 0;
			buffer[230] <= 0;
			buffer[231] <= 0;
			buffer[232] <= 0;
			buffer[233] <= 0;
			buffer[234] <= 0;
			buffer[235] <= 0;
			buffer[236] <= 0;
			buffer[237] <= 0;
			buffer[238] <= 0;
			buffer[239] <= 0;
			buffer[240] <= 0;
			buffer[241] <= 0;
			buffer[242] <= 0;
			buffer[243] <= 0;
			buffer[244] <= 0;
			buffer[245] <= 0;
			buffer[246] <= 0;
			buffer[247] <= 0;
			buffer[248] <= 0;
			buffer[249] <= 0;
			buffer[250] <= 0;
			buffer[251] <= 0;
			buffer[252] <= 0;
			buffer[253] <= 0;
			buffer[254] <= 0;
			buffer[255] <= 0;
			buffer[256] <= 0;
			buffer[257] <= 0;
			buffer[258] <= 0;
			buffer[259] <= 0;
			buffer[260] <= 0;
			buffer[261] <= 0;
			buffer[262] <= 0;
			buffer[263] <= 0;
			buffer[264] <= 0;
			buffer[265] <= 0;
			buffer[266] <= 0;
			buffer[267] <= 0;
			buffer[268] <= 0;
			buffer[269] <= 0;
			buffer[270] <= 0;
			buffer[271] <= 0;
			buffer[272] <= 0;
			buffer[273] <= 0;
			buffer[274] <= 0;
			buffer[275] <= 0;
			buffer[276] <= 0;
			buffer[277] <= 0;
			buffer[278] <= 0;
			buffer[279] <= 0;
			buffer[280] <= 0;
			buffer[281] <= 0;
			buffer[282] <= 0;
			buffer[283] <= 0;
			buffer[284] <= 0;
			buffer[285] <= 0;
			buffer[286] <= 0;
			buffer[287] <= 0;
		end else begin
			if (i_activation_in_en) begin
				buffer[i_counter * 4]     <= i_data[31:24];
				buffer[i_counter * 4 + 1] <= i_data[23:16];
				buffer[i_counter * 4 + 2] <= i_data[15:8];
				buffer[i_counter * 4 + 3] <= i_data[7:0];
			end
		end
	end

	
	wire [2:0] counter;
	assign counter = i_counter[5:3] - 1;

	always @(*) begin
		if (i_activation_out_en) begin
			if (counter == 3'd0) begin
				o_data = {buffer[  0][0],
					      buffer[  1][0],
						  buffer[  2][0],
						  buffer[  3][0],
						  buffer[  4][0],
						  buffer[  5][0],
						  buffer[  6][0],
						  buffer[  7][0],
						  buffer[  8][0],
						  buffer[  9][0],
						  buffer[ 10][0],
						  buffer[ 11][0],
						  buffer[ 12][0],
						  buffer[ 13][0],
						  buffer[ 14][0],
						  buffer[ 15][0],
						  buffer[ 16][0],
						  buffer[ 17][0],
						  buffer[ 18][0],
						  buffer[ 19][0],
						  buffer[ 20][0],
						  buffer[ 21][0],
						  buffer[ 22][0],
						  buffer[ 23][0],
						  buffer[ 24][0],
						  buffer[ 25][0],
						  buffer[ 26][0],
						  buffer[ 27][0],
						  buffer[ 28][0],
						  buffer[ 29][0],
						  buffer[ 30][0],
						  buffer[ 31][0],
						  buffer[ 32][0],
						  buffer[ 33][0],
						  buffer[ 34][0],
						  buffer[ 35][0],
						  buffer[ 36][0],
						  buffer[ 37][0],
						  buffer[ 38][0],
						  buffer[ 39][0],
						  buffer[ 40][0],
						  buffer[ 41][0],
						  buffer[ 42][0],
						  buffer[ 43][0],
						  buffer[ 44][0],
						  buffer[ 45][0],
						  buffer[ 46][0],
						  buffer[ 47][0],
						  buffer[ 48][0],
						  buffer[ 49][0],
						  buffer[ 50][0],
						  buffer[ 51][0],
						  buffer[ 52][0],
						  buffer[ 53][0],
						  buffer[ 54][0],
						  buffer[ 55][0],
						  buffer[ 56][0],
						  buffer[ 57][0],
						  buffer[ 58][0],
						  buffer[ 59][0],
						  buffer[ 60][0],
						  buffer[ 61][0],
						  buffer[ 62][0],
						  buffer[ 63][0],
						  buffer[ 64][0],
						  buffer[ 65][0],
						  buffer[ 66][0],
						  buffer[ 67][0],
						  buffer[ 68][0],
						  buffer[ 69][0],
						  buffer[ 70][0],
						  buffer[ 71][0],
						  buffer[ 72][0],
						  buffer[ 73][0],
						  buffer[ 74][0],
						  buffer[ 75][0],
						  buffer[ 76][0],
						  buffer[ 77][0],
						  buffer[ 78][0],
						  buffer[ 79][0],
						  buffer[ 80][0],
						  buffer[ 81][0],
						  buffer[ 82][0],
						  buffer[ 83][0],
						  buffer[ 84][0],
						  buffer[ 85][0],
						  buffer[ 86][0],
						  buffer[ 87][0],
						  buffer[ 88][0],
						  buffer[ 89][0],
						  buffer[ 90][0],
						  buffer[ 91][0],
						  buffer[ 92][0],
						  buffer[ 93][0],
						  buffer[ 94][0],
						  buffer[ 95][0],
						  buffer[ 96][0],
						  buffer[ 97][0],
						  buffer[ 98][0],
						  buffer[ 99][0],
						  buffer[100][0],
						  buffer[101][0],
						  buffer[102][0],
						  buffer[103][0],
						  buffer[104][0],
						  buffer[105][0],
						  buffer[106][0],
						  buffer[107][0],
						  buffer[108][0],
						  buffer[109][0],
						  buffer[110][0],
						  buffer[111][0],
						  buffer[112][0],
						  buffer[113][0],
						  buffer[114][0],
						  buffer[115][0],
						  buffer[116][0],
						  buffer[117][0],
						  buffer[118][0],
						  buffer[119][0],
						  buffer[120][0],
						  buffer[121][0],
						  buffer[122][0],
						  buffer[123][0],
						  buffer[124][0],
						  buffer[125][0],
						  buffer[126][0],
						  buffer[127][0],
						  buffer[128][0],
						  buffer[129][0],
						  buffer[130][0],
						  buffer[131][0],
						  buffer[132][0],
						  buffer[133][0],
						  buffer[134][0],
						  buffer[135][0],
						  buffer[136][0],
						  buffer[137][0],
						  buffer[138][0],
						  buffer[139][0],
						  buffer[140][0],
						  buffer[141][0],
						  buffer[142][0],
						  buffer[143][0],
						  buffer[144][0],
						  buffer[145][0],
						  buffer[146][0],
						  buffer[147][0],
						  buffer[148][0],
						  buffer[149][0],
						  buffer[150][0],
						  buffer[151][0],
						  buffer[152][0],
						  buffer[153][0],
						  buffer[154][0],
						  buffer[155][0],
						  buffer[156][0],
						  buffer[157][0],
						  buffer[158][0],
						  buffer[159][0],
						  buffer[160][0],
						  buffer[161][0],
						  buffer[162][0],
						  buffer[163][0],
						  buffer[164][0],
						  buffer[165][0],
						  buffer[166][0],
						  buffer[167][0],
						  buffer[168][0],
						  buffer[169][0],
						  buffer[170][0],
						  buffer[171][0],
						  buffer[172][0],
						  buffer[173][0],
						  buffer[174][0],
						  buffer[175][0],
						  buffer[176][0],
						  buffer[177][0],
						  buffer[178][0],
						  buffer[179][0],
						  buffer[180][0],
						  buffer[181][0],
						  buffer[182][0],
						  buffer[183][0],
						  buffer[184][0],
						  buffer[185][0],
						  buffer[186][0],
						  buffer[187][0],
						  buffer[188][0],
						  buffer[189][0],
						  buffer[190][0],
						  buffer[191][0],
						  buffer[192][0],
						  buffer[193][0],
						  buffer[194][0],
						  buffer[195][0],
						  buffer[196][0],
						  buffer[197][0],
						  buffer[198][0],
						  buffer[199][0],
						  buffer[200][0],
						  buffer[201][0],
						  buffer[202][0],
						  buffer[203][0],
						  buffer[204][0],
						  buffer[205][0],
						  buffer[206][0],
						  buffer[207][0],
						  buffer[208][0],
						  buffer[209][0],
						  buffer[210][0],
						  buffer[211][0],
						  buffer[212][0],
						  buffer[213][0],
						  buffer[214][0],
						  buffer[215][0],
						  buffer[216][0],
						  buffer[217][0],
						  buffer[218][0],
						  buffer[219][0],
						  buffer[220][0],
						  buffer[221][0],
						  buffer[222][0],
						  buffer[223][0],
						  buffer[224][0],
						  buffer[225][0],
						  buffer[226][0],
						  buffer[227][0],
						  buffer[228][0],
						  buffer[229][0],
						  buffer[230][0],
						  buffer[231][0],
						  buffer[232][0],
						  buffer[233][0],
						  buffer[234][0],
						  buffer[235][0],
						  buffer[236][0],
						  buffer[237][0],
						  buffer[238][0],
						  buffer[239][0],
						  buffer[240][0],
						  buffer[241][0],
						  buffer[242][0],
						  buffer[243][0],
						  buffer[244][0],
						  buffer[245][0],
						  buffer[246][0],
						  buffer[247][0],
						  buffer[248][0],
						  buffer[249][0],
						  buffer[250][0],
						  buffer[251][0],
						  buffer[252][0],
						  buffer[253][0],
						  buffer[254][0],
						  buffer[255][0],
						  buffer[256][0],
						  buffer[257][0],
						  buffer[258][0],
						  buffer[259][0],
						  buffer[260][0],
						  buffer[261][0],
						  buffer[262][0],
						  buffer[263][0],
						  buffer[264][0],
						  buffer[265][0],
						  buffer[266][0],
						  buffer[267][0],
						  buffer[268][0],
						  buffer[269][0],
						  buffer[270][0],
						  buffer[271][0],
						  buffer[272][0],
						  buffer[273][0],
						  buffer[274][0],
						  buffer[275][0],
						  buffer[276][0],
						  buffer[277][0],
						  buffer[278][0],
						  buffer[279][0],
						  buffer[280][0],
						  buffer[281][0],
						  buffer[282][0],
						  buffer[283][0],
						  buffer[284][0],
						  buffer[285][0],
						  buffer[286][0],
						  buffer[287][0]};
			end else if (counter == 3'd1) begin
				o_data = {buffer[  0][1],
					      buffer[  1][1],
						  buffer[  2][1],
						  buffer[  3][1],
						  buffer[  4][1],
						  buffer[  5][1],
						  buffer[  6][1],
						  buffer[  7][1],
						  buffer[  8][1],
						  buffer[  9][1],
						  buffer[ 10][1],
						  buffer[ 11][1],
						  buffer[ 12][1],
						  buffer[ 13][1],
						  buffer[ 14][1],
						  buffer[ 15][1],
						  buffer[ 16][1],
						  buffer[ 17][1],
						  buffer[ 18][1],
						  buffer[ 19][1],
						  buffer[ 20][1],
						  buffer[ 21][1],
						  buffer[ 22][1],
						  buffer[ 23][1],
						  buffer[ 24][1],
						  buffer[ 25][1],
						  buffer[ 26][1],
						  buffer[ 27][1],
						  buffer[ 28][1],
						  buffer[ 29][1],
						  buffer[ 30][1],
						  buffer[ 31][1],
						  buffer[ 32][1],
						  buffer[ 33][1],
						  buffer[ 34][1],
						  buffer[ 35][1],
						  buffer[ 36][1],
						  buffer[ 37][1],
						  buffer[ 38][1],
						  buffer[ 39][1],
						  buffer[ 40][1],
						  buffer[ 41][1],
						  buffer[ 42][1],
						  buffer[ 43][1],
						  buffer[ 44][1],
						  buffer[ 45][1],
						  buffer[ 46][1],
						  buffer[ 47][1],
						  buffer[ 48][1],
						  buffer[ 49][1],
						  buffer[ 50][1],
						  buffer[ 51][1],
						  buffer[ 52][1],
						  buffer[ 53][1],
						  buffer[ 54][1],
						  buffer[ 55][1],
						  buffer[ 56][1],
						  buffer[ 57][1],
						  buffer[ 58][1],
						  buffer[ 59][1],
						  buffer[ 60][1],
						  buffer[ 61][1],
						  buffer[ 62][1],
						  buffer[ 63][1],
						  buffer[ 64][1],
						  buffer[ 65][1],
						  buffer[ 66][1],
						  buffer[ 67][1],
						  buffer[ 68][1],
						  buffer[ 69][1],
						  buffer[ 70][1],
						  buffer[ 71][1],
						  buffer[ 72][1],
						  buffer[ 73][1],
						  buffer[ 74][1],
						  buffer[ 75][1],
						  buffer[ 76][1],
						  buffer[ 77][1],
						  buffer[ 78][1],
						  buffer[ 79][1],
						  buffer[ 80][1],
						  buffer[ 81][1],
						  buffer[ 82][1],
						  buffer[ 83][1],
						  buffer[ 84][1],
						  buffer[ 85][1],
						  buffer[ 86][1],
						  buffer[ 87][1],
						  buffer[ 88][1],
						  buffer[ 89][1],
						  buffer[ 90][1],
						  buffer[ 91][1],
						  buffer[ 92][1],
						  buffer[ 93][1],
						  buffer[ 94][1],
						  buffer[ 95][1],
						  buffer[ 96][1],
						  buffer[ 97][1],
						  buffer[ 98][1],
						  buffer[ 99][1],
						  buffer[100][1],
						  buffer[101][1],
						  buffer[102][1],
						  buffer[103][1],
						  buffer[104][1],
						  buffer[105][1],
						  buffer[106][1],
						  buffer[107][1],
						  buffer[108][1],
						  buffer[109][1],
						  buffer[110][1],
						  buffer[111][1],
						  buffer[112][1],
						  buffer[113][1],
						  buffer[114][1],
						  buffer[115][1],
						  buffer[116][1],
						  buffer[117][1],
						  buffer[118][1],
						  buffer[119][1],
						  buffer[120][1],
						  buffer[121][1],
						  buffer[122][1],
						  buffer[123][1],
						  buffer[124][1],
						  buffer[125][1],
						  buffer[126][1],
						  buffer[127][1],
						  buffer[128][1],
						  buffer[129][1],
						  buffer[130][1],
						  buffer[131][1],
						  buffer[132][1],
						  buffer[133][1],
						  buffer[134][1],
						  buffer[135][1],
						  buffer[136][1],
						  buffer[137][1],
						  buffer[138][1],
						  buffer[139][1],
						  buffer[140][1],
						  buffer[141][1],
						  buffer[142][1],
						  buffer[143][1],
						  buffer[144][1],
						  buffer[145][1],
						  buffer[146][1],
						  buffer[147][1],
						  buffer[148][1],
						  buffer[149][1],
						  buffer[150][1],
						  buffer[151][1],
						  buffer[152][1],
						  buffer[153][1],
						  buffer[154][1],
						  buffer[155][1],
						  buffer[156][1],
						  buffer[157][1],
						  buffer[158][1],
						  buffer[159][1],
						  buffer[160][1],
						  buffer[161][1],
						  buffer[162][1],
						  buffer[163][1],
						  buffer[164][1],
						  buffer[165][1],
						  buffer[166][1],
						  buffer[167][1],
						  buffer[168][1],
						  buffer[169][1],
						  buffer[170][1],
						  buffer[171][1],
						  buffer[172][1],
						  buffer[173][1],
						  buffer[174][1],
						  buffer[175][1],
						  buffer[176][1],
						  buffer[177][1],
						  buffer[178][1],
						  buffer[179][1],
						  buffer[180][1],
						  buffer[181][1],
						  buffer[182][1],
						  buffer[183][1],
						  buffer[184][1],
						  buffer[185][1],
						  buffer[186][1],
						  buffer[187][1],
						  buffer[188][1],
						  buffer[189][1],
						  buffer[190][1],
						  buffer[191][1],
						  buffer[192][1],
						  buffer[193][1],
						  buffer[194][1],
						  buffer[195][1],
						  buffer[196][1],
						  buffer[197][1],
						  buffer[198][1],
						  buffer[199][1],
						  buffer[200][1],
						  buffer[201][1],
						  buffer[202][1],
						  buffer[203][1],
						  buffer[204][1],
						  buffer[205][1],
						  buffer[206][1],
						  buffer[207][1],
						  buffer[208][1],
						  buffer[209][1],
						  buffer[210][1],
						  buffer[211][1],
						  buffer[212][1],
						  buffer[213][1],
						  buffer[214][1],
						  buffer[215][1],
						  buffer[216][1],
						  buffer[217][1],
						  buffer[218][1],
						  buffer[219][1],
						  buffer[220][1],
						  buffer[221][1],
						  buffer[222][1],
						  buffer[223][1],
						  buffer[224][1],
						  buffer[225][1],
						  buffer[226][1],
						  buffer[227][1],
						  buffer[228][1],
						  buffer[229][1],
						  buffer[230][1],
						  buffer[231][1],
						  buffer[232][1],
						  buffer[233][1],
						  buffer[234][1],
						  buffer[235][1],
						  buffer[236][1],
						  buffer[237][1],
						  buffer[238][1],
						  buffer[239][1],
						  buffer[240][1],
						  buffer[241][1],
						  buffer[242][1],
						  buffer[243][1],
						  buffer[244][1],
						  buffer[245][1],
						  buffer[246][1],
						  buffer[247][1],
						  buffer[248][1],
						  buffer[249][1],
						  buffer[250][1],
						  buffer[251][1],
						  buffer[252][1],
						  buffer[253][1],
						  buffer[254][1],
						  buffer[255][1],
						  buffer[256][1],
						  buffer[257][1],
						  buffer[258][1],
						  buffer[259][1],
						  buffer[260][1],
						  buffer[261][1],
						  buffer[262][1],
						  buffer[263][1],
						  buffer[264][1],
						  buffer[265][1],
						  buffer[266][1],
						  buffer[267][1],
						  buffer[268][1],
						  buffer[269][1],
						  buffer[270][1],
						  buffer[271][1],
						  buffer[272][1],
						  buffer[273][1],
						  buffer[274][1],
						  buffer[275][1],
						  buffer[276][1],
						  buffer[277][1],
						  buffer[278][1],
						  buffer[279][1],
						  buffer[280][1],
						  buffer[281][1],
						  buffer[282][1],
						  buffer[283][1],
						  buffer[284][1],
						  buffer[285][1],
						  buffer[286][1],
						  buffer[287][1]};
			end else if (counter == 3'd2) begin
				o_data = {buffer[  0][2],
					      buffer[  1][2],
						  buffer[  2][2],
						  buffer[  3][2],
						  buffer[  4][2],
						  buffer[  5][2],
						  buffer[  6][2],
						  buffer[  7][2],
						  buffer[  8][2],
						  buffer[  9][2],
						  buffer[ 10][2],
						  buffer[ 11][2],
						  buffer[ 12][2],
						  buffer[ 13][2],
						  buffer[ 14][2],
						  buffer[ 15][2],
						  buffer[ 16][2],
						  buffer[ 17][2],
						  buffer[ 18][2],
						  buffer[ 19][2],
						  buffer[ 20][2],
						  buffer[ 21][2],
						  buffer[ 22][2],
						  buffer[ 23][2],
						  buffer[ 24][2],
						  buffer[ 25][2],
						  buffer[ 26][2],
						  buffer[ 27][2],
						  buffer[ 28][2],
						  buffer[ 29][2],
						  buffer[ 30][2],
						  buffer[ 31][2],
						  buffer[ 32][2],
						  buffer[ 33][2],
						  buffer[ 34][2],
						  buffer[ 35][2],
						  buffer[ 36][2],
						  buffer[ 37][2],
						  buffer[ 38][2],
						  buffer[ 39][2],
						  buffer[ 40][2],
						  buffer[ 41][2],
						  buffer[ 42][2],
						  buffer[ 43][2],
						  buffer[ 44][2],
						  buffer[ 45][2],
						  buffer[ 46][2],
						  buffer[ 47][2],
						  buffer[ 48][2],
						  buffer[ 49][2],
						  buffer[ 50][2],
						  buffer[ 51][2],
						  buffer[ 52][2],
						  buffer[ 53][2],
						  buffer[ 54][2],
						  buffer[ 55][2],
						  buffer[ 56][2],
						  buffer[ 57][2],
						  buffer[ 58][2],
						  buffer[ 59][2],
						  buffer[ 60][2],
						  buffer[ 61][2],
						  buffer[ 62][2],
						  buffer[ 63][2],
						  buffer[ 64][2],
						  buffer[ 65][2],
						  buffer[ 66][2],
						  buffer[ 67][2],
						  buffer[ 68][2],
						  buffer[ 69][2],
						  buffer[ 70][2],
						  buffer[ 71][2],
						  buffer[ 72][2],
						  buffer[ 73][2],
						  buffer[ 74][2],
						  buffer[ 75][2],
						  buffer[ 76][2],
						  buffer[ 77][2],
						  buffer[ 78][2],
						  buffer[ 79][2],
						  buffer[ 80][2],
						  buffer[ 81][2],
						  buffer[ 82][2],
						  buffer[ 83][2],
						  buffer[ 84][2],
						  buffer[ 85][2],
						  buffer[ 86][2],
						  buffer[ 87][2],
						  buffer[ 88][2],
						  buffer[ 89][2],
						  buffer[ 90][2],
						  buffer[ 91][2],
						  buffer[ 92][2],
						  buffer[ 93][2],
						  buffer[ 94][2],
						  buffer[ 95][2],
						  buffer[ 96][2],
						  buffer[ 97][2],
						  buffer[ 98][2],
						  buffer[ 99][2],
						  buffer[100][2],
						  buffer[101][2],
						  buffer[102][2],
						  buffer[103][2],
						  buffer[104][2],
						  buffer[105][2],
						  buffer[106][2],
						  buffer[107][2],
						  buffer[108][2],
						  buffer[109][2],
						  buffer[110][2],
						  buffer[111][2],
						  buffer[112][2],
						  buffer[113][2],
						  buffer[114][2],
						  buffer[115][2],
						  buffer[116][2],
						  buffer[117][2],
						  buffer[118][2],
						  buffer[119][2],
						  buffer[120][2],
						  buffer[121][2],
						  buffer[122][2],
						  buffer[123][2],
						  buffer[124][2],
						  buffer[125][2],
						  buffer[126][2],
						  buffer[127][2],
						  buffer[128][2],
						  buffer[129][2],
						  buffer[130][2],
						  buffer[131][2],
						  buffer[132][2],
						  buffer[133][2],
						  buffer[134][2],
						  buffer[135][2],
						  buffer[136][2],
						  buffer[137][2],
						  buffer[138][2],
						  buffer[139][2],
						  buffer[140][2],
						  buffer[141][2],
						  buffer[142][2],
						  buffer[143][2],
						  buffer[144][2],
						  buffer[145][2],
						  buffer[146][2],
						  buffer[147][2],
						  buffer[148][2],
						  buffer[149][2],
						  buffer[150][2],
						  buffer[151][2],
						  buffer[152][2],
						  buffer[153][2],
						  buffer[154][2],
						  buffer[155][2],
						  buffer[156][2],
						  buffer[157][2],
						  buffer[158][2],
						  buffer[159][2],
						  buffer[160][2],
						  buffer[161][2],
						  buffer[162][2],
						  buffer[163][2],
						  buffer[164][2],
						  buffer[165][2],
						  buffer[166][2],
						  buffer[167][2],
						  buffer[168][2],
						  buffer[169][2],
						  buffer[170][2],
						  buffer[171][2],
						  buffer[172][2],
						  buffer[173][2],
						  buffer[174][2],
						  buffer[175][2],
						  buffer[176][2],
						  buffer[177][2],
						  buffer[178][2],
						  buffer[179][2],
						  buffer[180][2],
						  buffer[181][2],
						  buffer[182][2],
						  buffer[183][2],
						  buffer[184][2],
						  buffer[185][2],
						  buffer[186][2],
						  buffer[187][2],
						  buffer[188][2],
						  buffer[189][2],
						  buffer[190][2],
						  buffer[191][2],
						  buffer[192][2],
						  buffer[193][2],
						  buffer[194][2],
						  buffer[195][2],
						  buffer[196][2],
						  buffer[197][2],
						  buffer[198][2],
						  buffer[199][2],
						  buffer[200][2],
						  buffer[201][2],
						  buffer[202][2],
						  buffer[203][2],
						  buffer[204][2],
						  buffer[205][2],
						  buffer[206][2],
						  buffer[207][2],
						  buffer[208][2],
						  buffer[209][2],
						  buffer[210][2],
						  buffer[211][2],
						  buffer[212][2],
						  buffer[213][2],
						  buffer[214][2],
						  buffer[215][2],
						  buffer[216][2],
						  buffer[217][2],
						  buffer[218][2],
						  buffer[219][2],
						  buffer[220][2],
						  buffer[221][2],
						  buffer[222][2],
						  buffer[223][2],
						  buffer[224][2],
						  buffer[225][2],
						  buffer[226][2],
						  buffer[227][2],
						  buffer[228][2],
						  buffer[229][2],
						  buffer[230][2],
						  buffer[231][2],
						  buffer[232][2],
						  buffer[233][2],
						  buffer[234][2],
						  buffer[235][2],
						  buffer[236][2],
						  buffer[237][2],
						  buffer[238][2],
						  buffer[239][2],
						  buffer[240][2],
						  buffer[241][2],
						  buffer[242][2],
						  buffer[243][2],
						  buffer[244][2],
						  buffer[245][2],
						  buffer[246][2],
						  buffer[247][2],
						  buffer[248][2],
						  buffer[249][2],
						  buffer[250][2],
						  buffer[251][2],
						  buffer[252][2],
						  buffer[253][2],
						  buffer[254][2],
						  buffer[255][2],
						  buffer[256][2],
						  buffer[257][2],
						  buffer[258][2],
						  buffer[259][2],
						  buffer[260][2],
						  buffer[261][2],
						  buffer[262][2],
						  buffer[263][2],
						  buffer[264][2],
						  buffer[265][2],
						  buffer[266][2],
						  buffer[267][2],
						  buffer[268][2],
						  buffer[269][2],
						  buffer[270][2],
						  buffer[271][2],
						  buffer[272][2],
						  buffer[273][2],
						  buffer[274][2],
						  buffer[275][2],
						  buffer[276][2],
						  buffer[277][2],
						  buffer[278][2],
						  buffer[279][2],
						  buffer[280][2],
						  buffer[281][2],
						  buffer[282][2],
						  buffer[283][2],
						  buffer[284][2],
						  buffer[285][2],
						  buffer[286][2],
						  buffer[287][2]};
			end else if (counter == 3'd3) begin
				o_data = {buffer[  0][3],
					      buffer[  1][3],
						  buffer[  2][3],
						  buffer[  3][3],
						  buffer[  4][3],
						  buffer[  5][3],
						  buffer[  6][3],
						  buffer[  7][3],
						  buffer[  8][3],
						  buffer[  9][3],
						  buffer[ 10][3],
						  buffer[ 11][3],
						  buffer[ 12][3],
						  buffer[ 13][3],
						  buffer[ 14][3],
						  buffer[ 15][3],
						  buffer[ 16][3],
						  buffer[ 17][3],
						  buffer[ 18][3],
						  buffer[ 19][3],
						  buffer[ 20][3],
						  buffer[ 21][3],
						  buffer[ 22][3],
						  buffer[ 23][3],
						  buffer[ 24][3],
						  buffer[ 25][3],
						  buffer[ 26][3],
						  buffer[ 27][3],
						  buffer[ 28][3],
						  buffer[ 29][3],
						  buffer[ 30][3],
						  buffer[ 31][3],
						  buffer[ 32][3],
						  buffer[ 33][3],
						  buffer[ 34][3],
						  buffer[ 35][3],
						  buffer[ 36][3],
						  buffer[ 37][3],
						  buffer[ 38][3],
						  buffer[ 39][3],
						  buffer[ 40][3],
						  buffer[ 41][3],
						  buffer[ 42][3],
						  buffer[ 43][3],
						  buffer[ 44][3],
						  buffer[ 45][3],
						  buffer[ 46][3],
						  buffer[ 47][3],
						  buffer[ 48][3],
						  buffer[ 49][3],
						  buffer[ 50][3],
						  buffer[ 51][3],
						  buffer[ 52][3],
						  buffer[ 53][3],
						  buffer[ 54][3],
						  buffer[ 55][3],
						  buffer[ 56][3],
						  buffer[ 57][3],
						  buffer[ 58][3],
						  buffer[ 59][3],
						  buffer[ 60][3],
						  buffer[ 61][3],
						  buffer[ 62][3],
						  buffer[ 63][3],
						  buffer[ 64][3],
						  buffer[ 65][3],
						  buffer[ 66][3],
						  buffer[ 67][3],
						  buffer[ 68][3],
						  buffer[ 69][3],
						  buffer[ 70][3],
						  buffer[ 71][3],
						  buffer[ 72][3],
						  buffer[ 73][3],
						  buffer[ 74][3],
						  buffer[ 75][3],
						  buffer[ 76][3],
						  buffer[ 77][3],
						  buffer[ 78][3],
						  buffer[ 79][3],
						  buffer[ 80][3],
						  buffer[ 81][3],
						  buffer[ 82][3],
						  buffer[ 83][3],
						  buffer[ 84][3],
						  buffer[ 85][3],
						  buffer[ 86][3],
						  buffer[ 87][3],
						  buffer[ 88][3],
						  buffer[ 89][3],
						  buffer[ 90][3],
						  buffer[ 91][3],
						  buffer[ 92][3],
						  buffer[ 93][3],
						  buffer[ 94][3],
						  buffer[ 95][3],
						  buffer[ 96][3],
						  buffer[ 97][3],
						  buffer[ 98][3],
						  buffer[ 99][3],
						  buffer[100][3],
						  buffer[101][3],
						  buffer[102][3],
						  buffer[103][3],
						  buffer[104][3],
						  buffer[105][3],
						  buffer[106][3],
						  buffer[107][3],
						  buffer[108][3],
						  buffer[109][3],
						  buffer[110][3],
						  buffer[111][3],
						  buffer[112][3],
						  buffer[113][3],
						  buffer[114][3],
						  buffer[115][3],
						  buffer[116][3],
						  buffer[117][3],
						  buffer[118][3],
						  buffer[119][3],
						  buffer[120][3],
						  buffer[121][3],
						  buffer[122][3],
						  buffer[123][3],
						  buffer[124][3],
						  buffer[125][3],
						  buffer[126][3],
						  buffer[127][3],
						  buffer[128][3],
						  buffer[129][3],
						  buffer[130][3],
						  buffer[131][3],
						  buffer[132][3],
						  buffer[133][3],
						  buffer[134][3],
						  buffer[135][3],
						  buffer[136][3],
						  buffer[137][3],
						  buffer[138][3],
						  buffer[139][3],
						  buffer[140][3],
						  buffer[141][3],
						  buffer[142][3],
						  buffer[143][3],
						  buffer[144][3],
						  buffer[145][3],
						  buffer[146][3],
						  buffer[147][3],
						  buffer[148][3],
						  buffer[149][3],
						  buffer[150][3],
						  buffer[151][3],
						  buffer[152][3],
						  buffer[153][3],
						  buffer[154][3],
						  buffer[155][3],
						  buffer[156][3],
						  buffer[157][3],
						  buffer[158][3],
						  buffer[159][3],
						  buffer[160][3],
						  buffer[161][3],
						  buffer[162][3],
						  buffer[163][3],
						  buffer[164][3],
						  buffer[165][3],
						  buffer[166][3],
						  buffer[167][3],
						  buffer[168][3],
						  buffer[169][3],
						  buffer[170][3],
						  buffer[171][3],
						  buffer[172][3],
						  buffer[173][3],
						  buffer[174][3],
						  buffer[175][3],
						  buffer[176][3],
						  buffer[177][3],
						  buffer[178][3],
						  buffer[179][3],
						  buffer[180][3],
						  buffer[181][3],
						  buffer[182][3],
						  buffer[183][3],
						  buffer[184][3],
						  buffer[185][3],
						  buffer[186][3],
						  buffer[187][3],
						  buffer[188][3],
						  buffer[189][3],
						  buffer[190][3],
						  buffer[191][3],
						  buffer[192][3],
						  buffer[193][3],
						  buffer[194][3],
						  buffer[195][3],
						  buffer[196][3],
						  buffer[197][3],
						  buffer[198][3],
						  buffer[199][3],
						  buffer[200][3],
						  buffer[201][3],
						  buffer[202][3],
						  buffer[203][3],
						  buffer[204][3],
						  buffer[205][3],
						  buffer[206][3],
						  buffer[207][3],
						  buffer[208][3],
						  buffer[209][3],
						  buffer[210][3],
						  buffer[211][3],
						  buffer[212][3],
						  buffer[213][3],
						  buffer[214][3],
						  buffer[215][3],
						  buffer[216][3],
						  buffer[217][3],
						  buffer[218][3],
						  buffer[219][3],
						  buffer[220][3],
						  buffer[221][3],
						  buffer[222][3],
						  buffer[223][3],
						  buffer[224][3],
						  buffer[225][3],
						  buffer[226][3],
						  buffer[227][3],
						  buffer[228][3],
						  buffer[229][3],
						  buffer[230][3],
						  buffer[231][3],
						  buffer[232][3],
						  buffer[233][3],
						  buffer[234][3],
						  buffer[235][3],
						  buffer[236][3],
						  buffer[237][3],
						  buffer[238][3],
						  buffer[239][3],
						  buffer[240][3],
						  buffer[241][3],
						  buffer[242][3],
						  buffer[243][3],
						  buffer[244][3],
						  buffer[245][3],
						  buffer[246][3],
						  buffer[247][3],
						  buffer[248][3],
						  buffer[249][3],
						  buffer[250][3],
						  buffer[251][3],
						  buffer[252][3],
						  buffer[253][3],
						  buffer[254][3],
						  buffer[255][3],
						  buffer[256][3],
						  buffer[257][3],
						  buffer[258][3],
						  buffer[259][3],
						  buffer[260][3],
						  buffer[261][3],
						  buffer[262][3],
						  buffer[263][3],
						  buffer[264][3],
						  buffer[265][3],
						  buffer[266][3],
						  buffer[267][3],
						  buffer[268][3],
						  buffer[269][3],
						  buffer[270][3],
						  buffer[271][3],
						  buffer[272][3],
						  buffer[273][3],
						  buffer[274][3],
						  buffer[275][3],
						  buffer[276][3],
						  buffer[277][3],
						  buffer[278][3],
						  buffer[279][3],
						  buffer[280][3],
						  buffer[281][3],
						  buffer[282][3],
						  buffer[283][3],
						  buffer[284][3],
						  buffer[285][3],
						  buffer[286][3],
						  buffer[287][3]};
			end else if (counter == 3'd4) begin
				o_data = {buffer[  0][4],
					      buffer[  1][4],
						  buffer[  2][4],
						  buffer[  3][4],
						  buffer[  4][4],
						  buffer[  5][4],
						  buffer[  6][4],
						  buffer[  7][4],
						  buffer[  8][4],
						  buffer[  9][4],
						  buffer[ 10][4],
						  buffer[ 11][4],
						  buffer[ 12][4],
						  buffer[ 13][4],
						  buffer[ 14][4],
						  buffer[ 15][4],
						  buffer[ 16][4],
						  buffer[ 17][4],
						  buffer[ 18][4],
						  buffer[ 19][4],
						  buffer[ 20][4],
						  buffer[ 21][4],
						  buffer[ 22][4],
						  buffer[ 23][4],
						  buffer[ 24][4],
						  buffer[ 25][4],
						  buffer[ 26][4],
						  buffer[ 27][4],
						  buffer[ 28][4],
						  buffer[ 29][4],
						  buffer[ 30][4],
						  buffer[ 31][4],
						  buffer[ 32][4],
						  buffer[ 33][4],
						  buffer[ 34][4],
						  buffer[ 35][4],
						  buffer[ 36][4],
						  buffer[ 37][4],
						  buffer[ 38][4],
						  buffer[ 39][4],
						  buffer[ 40][4],
						  buffer[ 41][4],
						  buffer[ 42][4],
						  buffer[ 43][4],
						  buffer[ 44][4],
						  buffer[ 45][4],
						  buffer[ 46][4],
						  buffer[ 47][4],
						  buffer[ 48][4],
						  buffer[ 49][4],
						  buffer[ 50][4],
						  buffer[ 51][4],
						  buffer[ 52][4],
						  buffer[ 53][4],
						  buffer[ 54][4],
						  buffer[ 55][4],
						  buffer[ 56][4],
						  buffer[ 57][4],
						  buffer[ 58][4],
						  buffer[ 59][4],
						  buffer[ 60][4],
						  buffer[ 61][4],
						  buffer[ 62][4],
						  buffer[ 63][4],
						  buffer[ 64][4],
						  buffer[ 65][4],
						  buffer[ 66][4],
						  buffer[ 67][4],
						  buffer[ 68][4],
						  buffer[ 69][4],
						  buffer[ 70][4],
						  buffer[ 71][4],
						  buffer[ 72][4],
						  buffer[ 73][4],
						  buffer[ 74][4],
						  buffer[ 75][4],
						  buffer[ 76][4],
						  buffer[ 77][4],
						  buffer[ 78][4],
						  buffer[ 79][4],
						  buffer[ 80][4],
						  buffer[ 81][4],
						  buffer[ 82][4],
						  buffer[ 83][4],
						  buffer[ 84][4],
						  buffer[ 85][4],
						  buffer[ 86][4],
						  buffer[ 87][4],
						  buffer[ 88][4],
						  buffer[ 89][4],
						  buffer[ 90][4],
						  buffer[ 91][4],
						  buffer[ 92][4],
						  buffer[ 93][4],
						  buffer[ 94][4],
						  buffer[ 95][4],
						  buffer[ 96][4],
						  buffer[ 97][4],
						  buffer[ 98][4],
						  buffer[ 99][4],
						  buffer[100][4],
						  buffer[101][4],
						  buffer[102][4],
						  buffer[103][4],
						  buffer[104][4],
						  buffer[105][4],
						  buffer[106][4],
						  buffer[107][4],
						  buffer[108][4],
						  buffer[109][4],
						  buffer[110][4],
						  buffer[111][4],
						  buffer[112][4],
						  buffer[113][4],
						  buffer[114][4],
						  buffer[115][4],
						  buffer[116][4],
						  buffer[117][4],
						  buffer[118][4],
						  buffer[119][4],
						  buffer[120][4],
						  buffer[121][4],
						  buffer[122][4],
						  buffer[123][4],
						  buffer[124][4],
						  buffer[125][4],
						  buffer[126][4],
						  buffer[127][4],
						  buffer[128][4],
						  buffer[129][4],
						  buffer[130][4],
						  buffer[131][4],
						  buffer[132][4],
						  buffer[133][4],
						  buffer[134][4],
						  buffer[135][4],
						  buffer[136][4],
						  buffer[137][4],
						  buffer[138][4],
						  buffer[139][4],
						  buffer[140][4],
						  buffer[141][4],
						  buffer[142][4],
						  buffer[143][4],
						  buffer[144][4],
						  buffer[145][4],
						  buffer[146][4],
						  buffer[147][4],
						  buffer[148][4],
						  buffer[149][4],
						  buffer[150][4],
						  buffer[151][4],
						  buffer[152][4],
						  buffer[153][4],
						  buffer[154][4],
						  buffer[155][4],
						  buffer[156][4],
						  buffer[157][4],
						  buffer[158][4],
						  buffer[159][4],
						  buffer[160][4],
						  buffer[161][4],
						  buffer[162][4],
						  buffer[163][4],
						  buffer[164][4],
						  buffer[165][4],
						  buffer[166][4],
						  buffer[167][4],
						  buffer[168][4],
						  buffer[169][4],
						  buffer[170][4],
						  buffer[171][4],
						  buffer[172][4],
						  buffer[173][4],
						  buffer[174][4],
						  buffer[175][4],
						  buffer[176][4],
						  buffer[177][4],
						  buffer[178][4],
						  buffer[179][4],
						  buffer[180][4],
						  buffer[181][4],
						  buffer[182][4],
						  buffer[183][4],
						  buffer[184][4],
						  buffer[185][4],
						  buffer[186][4],
						  buffer[187][4],
						  buffer[188][4],
						  buffer[189][4],
						  buffer[190][4],
						  buffer[191][4],
						  buffer[192][4],
						  buffer[193][4],
						  buffer[194][4],
						  buffer[195][4],
						  buffer[196][4],
						  buffer[197][4],
						  buffer[198][4],
						  buffer[199][4],
						  buffer[200][4],
						  buffer[201][4],
						  buffer[202][4],
						  buffer[203][4],
						  buffer[204][4],
						  buffer[205][4],
						  buffer[206][4],
						  buffer[207][4],
						  buffer[208][4],
						  buffer[209][4],
						  buffer[210][4],
						  buffer[211][4],
						  buffer[212][4],
						  buffer[213][4],
						  buffer[214][4],
						  buffer[215][4],
						  buffer[216][4],
						  buffer[217][4],
						  buffer[218][4],
						  buffer[219][4],
						  buffer[220][4],
						  buffer[221][4],
						  buffer[222][4],
						  buffer[223][4],
						  buffer[224][4],
						  buffer[225][4],
						  buffer[226][4],
						  buffer[227][4],
						  buffer[228][4],
						  buffer[229][4],
						  buffer[230][4],
						  buffer[231][4],
						  buffer[232][4],
						  buffer[233][4],
						  buffer[234][4],
						  buffer[235][4],
						  buffer[236][4],
						  buffer[237][4],
						  buffer[238][4],
						  buffer[239][4],
						  buffer[240][4],
						  buffer[241][4],
						  buffer[242][4],
						  buffer[243][4],
						  buffer[244][4],
						  buffer[245][4],
						  buffer[246][4],
						  buffer[247][4],
						  buffer[248][4],
						  buffer[249][4],
						  buffer[250][4],
						  buffer[251][4],
						  buffer[252][4],
						  buffer[253][4],
						  buffer[254][4],
						  buffer[255][4],
						  buffer[256][4],
						  buffer[257][4],
						  buffer[258][4],
						  buffer[259][4],
						  buffer[260][4],
						  buffer[261][4],
						  buffer[262][4],
						  buffer[263][4],
						  buffer[264][4],
						  buffer[265][4],
						  buffer[266][4],
						  buffer[267][4],
						  buffer[268][4],
						  buffer[269][4],
						  buffer[270][4],
						  buffer[271][4],
						  buffer[272][4],
						  buffer[273][4],
						  buffer[274][4],
						  buffer[275][4],
						  buffer[276][4],
						  buffer[277][4],
						  buffer[278][4],
						  buffer[279][4],
						  buffer[280][4],
						  buffer[281][4],
						  buffer[282][4],
						  buffer[283][4],
						  buffer[284][4],
						  buffer[285][4],
						  buffer[286][4],
						  buffer[287][4]};
			end else if (counter == 3'd5) begin
				o_data = {buffer[  0][5],
					      buffer[  1][5],
						  buffer[  2][5],
						  buffer[  3][5],
						  buffer[  4][5],
						  buffer[  5][5],
						  buffer[  6][5],
						  buffer[  7][5],
						  buffer[  8][5],
						  buffer[  9][5],
						  buffer[ 10][5],
						  buffer[ 11][5],
						  buffer[ 12][5],
						  buffer[ 13][5],
						  buffer[ 14][5],
						  buffer[ 15][5],
						  buffer[ 16][5],
						  buffer[ 17][5],
						  buffer[ 18][5],
						  buffer[ 19][5],
						  buffer[ 20][5],
						  buffer[ 21][5],
						  buffer[ 22][5],
						  buffer[ 23][5],
						  buffer[ 24][5],
						  buffer[ 25][5],
						  buffer[ 26][5],
						  buffer[ 27][5],
						  buffer[ 28][5],
						  buffer[ 29][5],
						  buffer[ 30][5],
						  buffer[ 31][5],
						  buffer[ 32][5],
						  buffer[ 33][5],
						  buffer[ 34][5],
						  buffer[ 35][5],
						  buffer[ 36][5],
						  buffer[ 37][5],
						  buffer[ 38][5],
						  buffer[ 39][5],
						  buffer[ 40][5],
						  buffer[ 41][5],
						  buffer[ 42][5],
						  buffer[ 43][5],
						  buffer[ 44][5],
						  buffer[ 45][5],
						  buffer[ 46][5],
						  buffer[ 47][5],
						  buffer[ 48][5],
						  buffer[ 49][5],
						  buffer[ 50][5],
						  buffer[ 51][5],
						  buffer[ 52][5],
						  buffer[ 53][5],
						  buffer[ 54][5],
						  buffer[ 55][5],
						  buffer[ 56][5],
						  buffer[ 57][5],
						  buffer[ 58][5],
						  buffer[ 59][5],
						  buffer[ 60][5],
						  buffer[ 61][5],
						  buffer[ 62][5],
						  buffer[ 63][5],
						  buffer[ 64][5],
						  buffer[ 65][5],
						  buffer[ 66][5],
						  buffer[ 67][5],
						  buffer[ 68][5],
						  buffer[ 69][5],
						  buffer[ 70][5],
						  buffer[ 71][5],
						  buffer[ 72][5],
						  buffer[ 73][5],
						  buffer[ 74][5],
						  buffer[ 75][5],
						  buffer[ 76][5],
						  buffer[ 77][5],
						  buffer[ 78][5],
						  buffer[ 79][5],
						  buffer[ 80][5],
						  buffer[ 81][5],
						  buffer[ 82][5],
						  buffer[ 83][5],
						  buffer[ 84][5],
						  buffer[ 85][5],
						  buffer[ 86][5],
						  buffer[ 87][5],
						  buffer[ 88][5],
						  buffer[ 89][5],
						  buffer[ 90][5],
						  buffer[ 91][5],
						  buffer[ 92][5],
						  buffer[ 93][5],
						  buffer[ 94][5],
						  buffer[ 95][5],
						  buffer[ 96][5],
						  buffer[ 97][5],
						  buffer[ 98][5],
						  buffer[ 99][5],
						  buffer[100][5],
						  buffer[101][5],
						  buffer[102][5],
						  buffer[103][5],
						  buffer[104][5],
						  buffer[105][5],
						  buffer[106][5],
						  buffer[107][5],
						  buffer[108][5],
						  buffer[109][5],
						  buffer[110][5],
						  buffer[111][5],
						  buffer[112][5],
						  buffer[113][5],
						  buffer[114][5],
						  buffer[115][5],
						  buffer[116][5],
						  buffer[117][5],
						  buffer[118][5],
						  buffer[119][5],
						  buffer[120][5],
						  buffer[121][5],
						  buffer[122][5],
						  buffer[123][5],
						  buffer[124][5],
						  buffer[125][5],
						  buffer[126][5],
						  buffer[127][5],
						  buffer[128][5],
						  buffer[129][5],
						  buffer[130][5],
						  buffer[131][5],
						  buffer[132][5],
						  buffer[133][5],
						  buffer[134][5],
						  buffer[135][5],
						  buffer[136][5],
						  buffer[137][5],
						  buffer[138][5],
						  buffer[139][5],
						  buffer[140][5],
						  buffer[141][5],
						  buffer[142][5],
						  buffer[143][5],
						  buffer[144][5],
						  buffer[145][5],
						  buffer[146][5],
						  buffer[147][5],
						  buffer[148][5],
						  buffer[149][5],
						  buffer[150][5],
						  buffer[151][5],
						  buffer[152][5],
						  buffer[153][5],
						  buffer[154][5],
						  buffer[155][5],
						  buffer[156][5],
						  buffer[157][5],
						  buffer[158][5],
						  buffer[159][5],
						  buffer[160][5],
						  buffer[161][5],
						  buffer[162][5],
						  buffer[163][5],
						  buffer[164][5],
						  buffer[165][5],
						  buffer[166][5],
						  buffer[167][5],
						  buffer[168][5],
						  buffer[169][5],
						  buffer[170][5],
						  buffer[171][5],
						  buffer[172][5],
						  buffer[173][5],
						  buffer[174][5],
						  buffer[175][5],
						  buffer[176][5],
						  buffer[177][5],
						  buffer[178][5],
						  buffer[179][5],
						  buffer[180][5],
						  buffer[181][5],
						  buffer[182][5],
						  buffer[183][5],
						  buffer[184][5],
						  buffer[185][5],
						  buffer[186][5],
						  buffer[187][5],
						  buffer[188][5],
						  buffer[189][5],
						  buffer[190][5],
						  buffer[191][5],
						  buffer[192][5],
						  buffer[193][5],
						  buffer[194][5],
						  buffer[195][5],
						  buffer[196][5],
						  buffer[197][5],
						  buffer[198][5],
						  buffer[199][5],
						  buffer[200][5],
						  buffer[201][5],
						  buffer[202][5],
						  buffer[203][5],
						  buffer[204][5],
						  buffer[205][5],
						  buffer[206][5],
						  buffer[207][5],
						  buffer[208][5],
						  buffer[209][5],
						  buffer[210][5],
						  buffer[211][5],
						  buffer[212][5],
						  buffer[213][5],
						  buffer[214][5],
						  buffer[215][5],
						  buffer[216][5],
						  buffer[217][5],
						  buffer[218][5],
						  buffer[219][5],
						  buffer[220][5],
						  buffer[221][5],
						  buffer[222][5],
						  buffer[223][5],
						  buffer[224][5],
						  buffer[225][5],
						  buffer[226][5],
						  buffer[227][5],
						  buffer[228][5],
						  buffer[229][5],
						  buffer[230][5],
						  buffer[231][5],
						  buffer[232][5],
						  buffer[233][5],
						  buffer[234][5],
						  buffer[235][5],
						  buffer[236][5],
						  buffer[237][5],
						  buffer[238][5],
						  buffer[239][5],
						  buffer[240][5],
						  buffer[241][5],
						  buffer[242][5],
						  buffer[243][5],
						  buffer[244][5],
						  buffer[245][5],
						  buffer[246][5],
						  buffer[247][5],
						  buffer[248][5],
						  buffer[249][5],
						  buffer[250][5],
						  buffer[251][5],
						  buffer[252][5],
						  buffer[253][5],
						  buffer[254][5],
						  buffer[255][5],
						  buffer[256][5],
						  buffer[257][5],
						  buffer[258][5],
						  buffer[259][5],
						  buffer[260][5],
						  buffer[261][5],
						  buffer[262][5],
						  buffer[263][5],
						  buffer[264][5],
						  buffer[265][5],
						  buffer[266][5],
						  buffer[267][5],
						  buffer[268][5],
						  buffer[269][5],
						  buffer[270][5],
						  buffer[271][5],
						  buffer[272][5],
						  buffer[273][5],
						  buffer[274][5],
						  buffer[275][5],
						  buffer[276][5],
						  buffer[277][5],
						  buffer[278][5],
						  buffer[279][5],
						  buffer[280][5],
						  buffer[281][5],
						  buffer[282][5],
						  buffer[283][5],
						  buffer[284][5],
						  buffer[285][5],
						  buffer[286][5],
						  buffer[287][5]};
			end else if (counter == 3'd6) begin
				o_data = {buffer[  0][6],
					      buffer[  1][6],
						  buffer[  2][6],
						  buffer[  3][6],
						  buffer[  4][6],
						  buffer[  5][6],
						  buffer[  6][6],
						  buffer[  7][6],
						  buffer[  8][6],
						  buffer[  9][6],
						  buffer[ 10][6],
						  buffer[ 11][6],
						  buffer[ 12][6],
						  buffer[ 13][6],
						  buffer[ 14][6],
						  buffer[ 15][6],
						  buffer[ 16][6],
						  buffer[ 17][6],
						  buffer[ 18][6],
						  buffer[ 19][6],
						  buffer[ 20][6],
						  buffer[ 21][6],
						  buffer[ 22][6],
						  buffer[ 23][6],
						  buffer[ 24][6],
						  buffer[ 25][6],
						  buffer[ 26][6],
						  buffer[ 27][6],
						  buffer[ 28][6],
						  buffer[ 29][6],
						  buffer[ 30][6],
						  buffer[ 31][6],
						  buffer[ 32][6],
						  buffer[ 33][6],
						  buffer[ 34][6],
						  buffer[ 35][6],
						  buffer[ 36][6],
						  buffer[ 37][6],
						  buffer[ 38][6],
						  buffer[ 39][6],
						  buffer[ 40][6],
						  buffer[ 41][6],
						  buffer[ 42][6],
						  buffer[ 43][6],
						  buffer[ 44][6],
						  buffer[ 45][6],
						  buffer[ 46][6],
						  buffer[ 47][6],
						  buffer[ 48][6],
						  buffer[ 49][6],
						  buffer[ 50][6],
						  buffer[ 51][6],
						  buffer[ 52][6],
						  buffer[ 53][6],
						  buffer[ 54][6],
						  buffer[ 55][6],
						  buffer[ 56][6],
						  buffer[ 57][6],
						  buffer[ 58][6],
						  buffer[ 59][6],
						  buffer[ 60][6],
						  buffer[ 61][6],
						  buffer[ 62][6],
						  buffer[ 63][6],
						  buffer[ 64][6],
						  buffer[ 65][6],
						  buffer[ 66][6],
						  buffer[ 67][6],
						  buffer[ 68][6],
						  buffer[ 69][6],
						  buffer[ 70][6],
						  buffer[ 71][6],
						  buffer[ 72][6],
						  buffer[ 73][6],
						  buffer[ 74][6],
						  buffer[ 75][6],
						  buffer[ 76][6],
						  buffer[ 77][6],
						  buffer[ 78][6],
						  buffer[ 79][6],
						  buffer[ 80][6],
						  buffer[ 81][6],
						  buffer[ 82][6],
						  buffer[ 83][6],
						  buffer[ 84][6],
						  buffer[ 85][6],
						  buffer[ 86][6],
						  buffer[ 87][6],
						  buffer[ 88][6],
						  buffer[ 89][6],
						  buffer[ 90][6],
						  buffer[ 91][6],
						  buffer[ 92][6],
						  buffer[ 93][6],
						  buffer[ 94][6],
						  buffer[ 95][6],
						  buffer[ 96][6],
						  buffer[ 97][6],
						  buffer[ 98][6],
						  buffer[ 99][6],
						  buffer[100][6],
						  buffer[101][6],
						  buffer[102][6],
						  buffer[103][6],
						  buffer[104][6],
						  buffer[105][6],
						  buffer[106][6],
						  buffer[107][6],
						  buffer[108][6],
						  buffer[109][6],
						  buffer[110][6],
						  buffer[111][6],
						  buffer[112][6],
						  buffer[113][6],
						  buffer[114][6],
						  buffer[115][6],
						  buffer[116][6],
						  buffer[117][6],
						  buffer[118][6],
						  buffer[119][6],
						  buffer[120][6],
						  buffer[121][6],
						  buffer[122][6],
						  buffer[123][6],
						  buffer[124][6],
						  buffer[125][6],
						  buffer[126][6],
						  buffer[127][6],
						  buffer[128][6],
						  buffer[129][6],
						  buffer[130][6],
						  buffer[131][6],
						  buffer[132][6],
						  buffer[133][6],
						  buffer[134][6],
						  buffer[135][6],
						  buffer[136][6],
						  buffer[137][6],
						  buffer[138][6],
						  buffer[139][6],
						  buffer[140][6],
						  buffer[141][6],
						  buffer[142][6],
						  buffer[143][6],
						  buffer[144][6],
						  buffer[145][6],
						  buffer[146][6],
						  buffer[147][6],
						  buffer[148][6],
						  buffer[149][6],
						  buffer[150][6],
						  buffer[151][6],
						  buffer[152][6],
						  buffer[153][6],
						  buffer[154][6],
						  buffer[155][6],
						  buffer[156][6],
						  buffer[157][6],
						  buffer[158][6],
						  buffer[159][6],
						  buffer[160][6],
						  buffer[161][6],
						  buffer[162][6],
						  buffer[163][6],
						  buffer[164][6],
						  buffer[165][6],
						  buffer[166][6],
						  buffer[167][6],
						  buffer[168][6],
						  buffer[169][6],
						  buffer[170][6],
						  buffer[171][6],
						  buffer[172][6],
						  buffer[173][6],
						  buffer[174][6],
						  buffer[175][6],
						  buffer[176][6],
						  buffer[177][6],
						  buffer[178][6],
						  buffer[179][6],
						  buffer[180][6],
						  buffer[181][6],
						  buffer[182][6],
						  buffer[183][6],
						  buffer[184][6],
						  buffer[185][6],
						  buffer[186][6],
						  buffer[187][6],
						  buffer[188][6],
						  buffer[189][6],
						  buffer[190][6],
						  buffer[191][6],
						  buffer[192][6],
						  buffer[193][6],
						  buffer[194][6],
						  buffer[195][6],
						  buffer[196][6],
						  buffer[197][6],
						  buffer[198][6],
						  buffer[199][6],
						  buffer[200][6],
						  buffer[201][6],
						  buffer[202][6],
						  buffer[203][6],
						  buffer[204][6],
						  buffer[205][6],
						  buffer[206][6],
						  buffer[207][6],
						  buffer[208][6],
						  buffer[209][6],
						  buffer[210][6],
						  buffer[211][6],
						  buffer[212][6],
						  buffer[213][6],
						  buffer[214][6],
						  buffer[215][6],
						  buffer[216][6],
						  buffer[217][6],
						  buffer[218][6],
						  buffer[219][6],
						  buffer[220][6],
						  buffer[221][6],
						  buffer[222][6],
						  buffer[223][6],
						  buffer[224][6],
						  buffer[225][6],
						  buffer[226][6],
						  buffer[227][6],
						  buffer[228][6],
						  buffer[229][6],
						  buffer[230][6],
						  buffer[231][6],
						  buffer[232][6],
						  buffer[233][6],
						  buffer[234][6],
						  buffer[235][6],
						  buffer[236][6],
						  buffer[237][6],
						  buffer[238][6],
						  buffer[239][6],
						  buffer[240][6],
						  buffer[241][6],
						  buffer[242][6],
						  buffer[243][6],
						  buffer[244][6],
						  buffer[245][6],
						  buffer[246][6],
						  buffer[247][6],
						  buffer[248][6],
						  buffer[249][6],
						  buffer[250][6],
						  buffer[251][6],
						  buffer[252][6],
						  buffer[253][6],
						  buffer[254][6],
						  buffer[255][6],
						  buffer[256][6],
						  buffer[257][6],
						  buffer[258][6],
						  buffer[259][6],
						  buffer[260][6],
						  buffer[261][6],
						  buffer[262][6],
						  buffer[263][6],
						  buffer[264][6],
						  buffer[265][6],
						  buffer[266][6],
						  buffer[267][6],
						  buffer[268][6],
						  buffer[269][6],
						  buffer[270][6],
						  buffer[271][6],
						  buffer[272][6],
						  buffer[273][6],
						  buffer[274][6],
						  buffer[275][6],
						  buffer[276][6],
						  buffer[277][6],
						  buffer[278][6],
						  buffer[279][6],
						  buffer[280][6],
						  buffer[281][6],
						  buffer[282][6],
						  buffer[283][6],
						  buffer[284][6],
						  buffer[285][6],
						  buffer[286][6],
						  buffer[287][6]};
			end else if (counter == 3'd7) begin
				o_data = {buffer[  0][7],
					      buffer[  1][7],
						  buffer[  2][7],
						  buffer[  3][7],
						  buffer[  4][7],
						  buffer[  5][7],
						  buffer[  6][7],
						  buffer[  7][7],
						  buffer[  8][7],
						  buffer[  9][7],
						  buffer[ 10][7],
						  buffer[ 11][7],
						  buffer[ 12][7],
						  buffer[ 13][7],
						  buffer[ 14][7],
						  buffer[ 15][7],
						  buffer[ 16][7],
						  buffer[ 17][7],
						  buffer[ 18][7],
						  buffer[ 19][7],
						  buffer[ 20][7],
						  buffer[ 21][7],
						  buffer[ 22][7],
						  buffer[ 23][7],
						  buffer[ 24][7],
						  buffer[ 25][7],
						  buffer[ 26][7],
						  buffer[ 27][7],
						  buffer[ 28][7],
						  buffer[ 29][7],
						  buffer[ 30][7],
						  buffer[ 31][7],
						  buffer[ 32][7],
						  buffer[ 33][7],
						  buffer[ 34][7],
						  buffer[ 35][7],
						  buffer[ 36][7],
						  buffer[ 37][7],
						  buffer[ 38][7],
						  buffer[ 39][7],
						  buffer[ 40][7],
						  buffer[ 41][7],
						  buffer[ 42][7],
						  buffer[ 43][7],
						  buffer[ 44][7],
						  buffer[ 45][7],
						  buffer[ 46][7],
						  buffer[ 47][7],
						  buffer[ 48][7],
						  buffer[ 49][7],
						  buffer[ 50][7],
						  buffer[ 51][7],
						  buffer[ 52][7],
						  buffer[ 53][7],
						  buffer[ 54][7],
						  buffer[ 55][7],
						  buffer[ 56][7],
						  buffer[ 57][7],
						  buffer[ 58][7],
						  buffer[ 59][7],
						  buffer[ 60][7],
						  buffer[ 61][7],
						  buffer[ 62][7],
						  buffer[ 63][7],
						  buffer[ 64][7],
						  buffer[ 65][7],
						  buffer[ 66][7],
						  buffer[ 67][7],
						  buffer[ 68][7],
						  buffer[ 69][7],
						  buffer[ 70][7],
						  buffer[ 71][7],
						  buffer[ 72][7],
						  buffer[ 73][7],
						  buffer[ 74][7],
						  buffer[ 75][7],
						  buffer[ 76][7],
						  buffer[ 77][7],
						  buffer[ 78][7],
						  buffer[ 79][7],
						  buffer[ 80][7],
						  buffer[ 81][7],
						  buffer[ 82][7],
						  buffer[ 83][7],
						  buffer[ 84][7],
						  buffer[ 85][7],
						  buffer[ 86][7],
						  buffer[ 87][7],
						  buffer[ 88][7],
						  buffer[ 89][7],
						  buffer[ 90][7],
						  buffer[ 91][7],
						  buffer[ 92][7],
						  buffer[ 93][7],
						  buffer[ 94][7],
						  buffer[ 95][7],
						  buffer[ 96][7],
						  buffer[ 97][7],
						  buffer[ 98][7],
						  buffer[ 99][7],
						  buffer[100][7],
						  buffer[101][7],
						  buffer[102][7],
						  buffer[103][7],
						  buffer[104][7],
						  buffer[105][7],
						  buffer[106][7],
						  buffer[107][7],
						  buffer[108][7],
						  buffer[109][7],
						  buffer[110][7],
						  buffer[111][7],
						  buffer[112][7],
						  buffer[113][7],
						  buffer[114][7],
						  buffer[115][7],
						  buffer[116][7],
						  buffer[117][7],
						  buffer[118][7],
						  buffer[119][7],
						  buffer[120][7],
						  buffer[121][7],
						  buffer[122][7],
						  buffer[123][7],
						  buffer[124][7],
						  buffer[125][7],
						  buffer[126][7],
						  buffer[127][7],
						  buffer[128][7],
						  buffer[129][7],
						  buffer[130][7],
						  buffer[131][7],
						  buffer[132][7],
						  buffer[133][7],
						  buffer[134][7],
						  buffer[135][7],
						  buffer[136][7],
						  buffer[137][7],
						  buffer[138][7],
						  buffer[139][7],
						  buffer[140][7],
						  buffer[141][7],
						  buffer[142][7],
						  buffer[143][7],
						  buffer[144][7],
						  buffer[145][7],
						  buffer[146][7],
						  buffer[147][7],
						  buffer[148][7],
						  buffer[149][7],
						  buffer[150][7],
						  buffer[151][7],
						  buffer[152][7],
						  buffer[153][7],
						  buffer[154][7],
						  buffer[155][7],
						  buffer[156][7],
						  buffer[157][7],
						  buffer[158][7],
						  buffer[159][7],
						  buffer[160][7],
						  buffer[161][7],
						  buffer[162][7],
						  buffer[163][7],
						  buffer[164][7],
						  buffer[165][7],
						  buffer[166][7],
						  buffer[167][7],
						  buffer[168][7],
						  buffer[169][7],
						  buffer[170][7],
						  buffer[171][7],
						  buffer[172][7],
						  buffer[173][7],
						  buffer[174][7],
						  buffer[175][7],
						  buffer[176][7],
						  buffer[177][7],
						  buffer[178][7],
						  buffer[179][7],
						  buffer[180][7],
						  buffer[181][7],
						  buffer[182][7],
						  buffer[183][7],
						  buffer[184][7],
						  buffer[185][7],
						  buffer[186][7],
						  buffer[187][7],
						  buffer[188][7],
						  buffer[189][7],
						  buffer[190][7],
						  buffer[191][7],
						  buffer[192][7],
						  buffer[193][7],
						  buffer[194][7],
						  buffer[195][7],
						  buffer[196][7],
						  buffer[197][7],
						  buffer[198][7],
						  buffer[199][7],
						  buffer[200][7],
						  buffer[201][7],
						  buffer[202][7],
						  buffer[203][7],
						  buffer[204][7],
						  buffer[205][7],
						  buffer[206][7],
						  buffer[207][7],
						  buffer[208][7],
						  buffer[209][7],
						  buffer[210][7],
						  buffer[211][7],
						  buffer[212][7],
						  buffer[213][7],
						  buffer[214][7],
						  buffer[215][7],
						  buffer[216][7],
						  buffer[217][7],
						  buffer[218][7],
						  buffer[219][7],
						  buffer[220][7],
						  buffer[221][7],
						  buffer[222][7],
						  buffer[223][7],
						  buffer[224][7],
						  buffer[225][7],
						  buffer[226][7],
						  buffer[227][7],
						  buffer[228][7],
						  buffer[229][7],
						  buffer[230][7],
						  buffer[231][7],
						  buffer[232][7],
						  buffer[233][7],
						  buffer[234][7],
						  buffer[235][7],
						  buffer[236][7],
						  buffer[237][7],
						  buffer[238][7],
						  buffer[239][7],
						  buffer[240][7],
						  buffer[241][7],
						  buffer[242][7],
						  buffer[243][7],
						  buffer[244][7],
						  buffer[245][7],
						  buffer[246][7],
						  buffer[247][7],
						  buffer[248][7],
						  buffer[249][7],
						  buffer[250][7],
						  buffer[251][7],
						  buffer[252][7],
						  buffer[253][7],
						  buffer[254][7],
						  buffer[255][7],
						  buffer[256][7],
						  buffer[257][7],
						  buffer[258][7],
						  buffer[259][7],
						  buffer[260][7],
						  buffer[261][7],
						  buffer[262][7],
						  buffer[263][7],
						  buffer[264][7],
						  buffer[265][7],
						  buffer[266][7],
						  buffer[267][7],
						  buffer[268][7],
						  buffer[269][7],
						  buffer[270][7],
						  buffer[271][7],
						  buffer[272][7],
						  buffer[273][7],
						  buffer[274][7],
						  buffer[275][7],
						  buffer[276][7],
						  buffer[277][7],
						  buffer[278][7],
						  buffer[279][7],
						  buffer[280][7],
						  buffer[281][7],
						  buffer[282][7],
						  buffer[283][7],
						  buffer[284][7],
						  buffer[285][7],
						  buffer[286][7],
						  buffer[287][7]};
			end
		end else begin
			o_data = 0;
		end
	end

endmodule






























/*
module activation_buffer (
	input i_clk,
	input i_rst,
	input i_activation_en,
	input [6:0] i_counter,
	input [31:0] i_data,
	output [287:0] o_data
);

	reg [7:0] buffer [0:287];

	always @(posedge i_clk) begin
		if (rst) begin
			buffer[0] <= 0;
			buffer[1] <= 0;
			buffer[2] <= 0;
			buffer[3] <= 0;
			buffer[4] <= 0;
			buffer[5] <= 0;
			buffer[6] <= 0;
			buffer[7] <= 0;
		end else begin
			if (i_activation_en) begin
				if (i_counter == 7'd0) begin
					buffer[0][287:284] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][287:284] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][287:284] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][287:284] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][287:284] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][287:284] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][287:284] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][287:284] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd1) begin
					buffer[0][283:280] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][283:280] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][283:280] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][283:280] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][283:280] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][283:280] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][283:280] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][283:280] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd2) begin
					buffer[0][279:276] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][279:276] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][279:276] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][279:276] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][279:276] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][279:276] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][279:276] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][279:276] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd3) begin
					buffer[0][275:272] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][275:272] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][275:272] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][275:272] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][275:272] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][275:272] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][275:272] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][275:272] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd4) begin
					buffer[0][271:268] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][271:268] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][271:268] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][271:268] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][271:268] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][271:268] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][271:268] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][271:268] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd5) begin
					buffer[0][267:264] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][267:264] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][267:264] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][267:264] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][267:264] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][267:264] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][267:264] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][267:264] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd6) begin
					buffer[0][263:260] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][263:260] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][263:260] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][263:260] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][263:260] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][263:260] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][263:260] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][263:260] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd7) begin
					buffer[0][259:256] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][259:256] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][259:256] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][259:256] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][259:256] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][259:256] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][259:256] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][259:256] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd8) begin
					buffer[0][255:252] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][255:252] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][255:252] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][255:252] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][255:252] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][255:252] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][255:252] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][255:252] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd9) begin
					buffer[0][251:248] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][251:248] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][251:248] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][251:248] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][251:248] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][251:248] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][251:248] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][251:248] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd10) begin
					buffer[0][247:244] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][247:244] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][247:244] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][247:244] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][247:244] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][247:244] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][247:244] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][247:244] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd11) begin
					buffer[0][243:240] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][243:240] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][243:240] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][243:240] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][243:240] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][243:240] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][243:240] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][243:240] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd12) begin
					buffer[0][239:236] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][239:236] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][239:236] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][239:236] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][239:236] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][239:236] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][239:236] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][239:236] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd13) begin
					buffer[0][235:232] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][235:232] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][235:232] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][235:232] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][235:232] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][235:232] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][235:232] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][235:232] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd14) begin
					buffer[0][231:228] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][231:228] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][231:228] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][231:228] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][231:228] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][231:228] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][231:228] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][231:228] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd14) begin
					buffer[0][231:228] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][231:228] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][231:228] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][231:228] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][231:228] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][231:228] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][231:228] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][231:228] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd15) begin
					buffer[0][237:224] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][237:224] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][237:224] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][237:224] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][237:224] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][237:224] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][237:224] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][237:224] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end else if (i_counter == 7'd16) begin
					buffer[0][237:223] <= {i_data[24], i_data[16], i_data[8],  i_data[0]};
					buffer[1][237:223] <= {i_data[25], i_data[17], i_data[9],  i_data[1]};
					buffer[2][237:223] <= {i_data[26], i_data[18], i_data[10], i_data[2]};
					buffer[3][237:223] <= {i_data[27], i_data[19], i_data[11], i_data[3]};
					buffer[4][237:223] <= {i_data[28], i_data[20], i_data[12], i_data[4]};
					buffer[5][237:223] <= {i_data[29], i_data[21], i_data[13], i_data[5]};
					buffer[6][237:223] <= {i_data[30], i_data[22], i_data[14], i_data[6]};
					buffer[7][237:223] <= {i_data[31], i_data[23], i_data[15], i_data[7]};
				end
			end
		end
	end
	assign o_data = (i_compute_en && i_counter[2:0] == 3'b111) ? buffer[i_counter[5:3]] : 288'b0


endmodule

*/

