module PIM_TOP (
	input i_clk, 
	input i_rst,

	//RISCV I/O
	input [31:0] i_address,
	input [31:0] i_data,
	output [31:0] o_data,

	//weight
	output o_weight_out_en0,
	output o_weight_out_en1,
	output o_weight_out_en2,
	output o_weight_out_en3,
	output [8:0] o_WL_address0,
	output [8:0] o_WL_address1,
	output [8:0] o_WL_address2,
	output [8:0] o_WL_address3,
	output [255:0] o_cam_data0,
	output [255:0] o_cam_data1,
	output [255:0] o_cam_data2,
	output [255:0] o_cam_data3,
	output [255:0] o_cim_data0,
	output [255:0] o_cim_data1,
	output [255:0] o_cim_data2,
	output [255:0] o_cim_data3,

	//activation
	output o_activation_out_en0,
	output o_activation_out_en1,
	output o_activation_out_en2,
	output o_activation_out_en3,
	output [287:0] o_activation_out_data0,
	output [287:0] o_activation_out_data1,
	output [287:0] o_activation_out_data2,
	output [287:0] o_activation_out_data3,

	//result
	input [31:0] result0,
	input [31:0] result1,
	input [31:0] result2,
	input [31:0] result3,
	input [31:0] result4,
	input [31:0] result5,
	input [31:0] result6,
	input [31:0] result7,
	input [31:0] result8,
	input [31:0] result9,
	input [31:0] result10,
	input [31:0] result11,
	input [31:0] result12,
	input [31:0] result13,
	input [31:0] result14,
	input [31:0] result15,
	input [31:0] result16,
	input [31:0] result17,
	input [31:0] result18,
	input [31:0] result19,
	input [31:0] result20,
	input [31:0] result21,
	input [31:0] result22,
	input [31:0] result23,
	input [31:0] result24,
	input [31:0] result25,
	input [31:0] result26,
	input [31:0] result27,
	input [31:0] result28,
	input [31:0] result29,
	input [31:0] result30,
	input [31:0] result31,
	input [31:0] result32,
	input [31:0] result33,
	input [31:0] result34,
	input [31:0] result35,
	input [31:0] result36,
	input [31:0] result37,
	input [31:0] result38,
	input [31:0] result39,
	input [31:0] result40,
	input [31:0] result41,
	input [31:0] result42,
	input [31:0] result43,
	input [31:0] result44,
	input [31:0] result45,
	input [31:0] result46,
	input [31:0] result47,
	input [31:0] result48,
	input [31:0] result49,
	input [31:0] result50,
	input [31:0] result51,
	input [31:0] result52,
	input [31:0] result53,
	input [31:0] result54,
	input [31:0] result55,
	input [31:0] result56,
	input [31:0] result57,
	input [31:0] result58,
	input [31:0] result59,
	input [31:0] result60,
	input [31:0] result61,
	input [31:0] result62,
	input [31:0] result63,
	input [31:0] result64,
	input [31:0] result65,
	input [31:0] result66,
	input [31:0] result67,
	input [31:0] result68,
	input [31:0] result69,
	input [31:0] result70,
	input [31:0] result71,
	input [31:0] result72,
	input [31:0] result73,
	input [31:0] result74,
	input [31:0] result75,
	input [31:0] result76,
	input [31:0] result77,
	input [31:0] result78,
	input [31:0] result79,
	input [31:0] result80,
	input [31:0] result81,
	input [31:0] result82,
	input [31:0] result83,
	input [31:0] result84,
	input [31:0] result85,
	input [31:0] result86,
	input [31:0] result87,
	input [31:0] result88,
	input [31:0] result89,
	input [31:0] result90,
	input [31:0] result91,
	input [31:0] result92,
	input [31:0] result93,
	input [31:0] result94,
	input [31:0] result95,
	input [31:0] result96,
	input [31:0] result97,
	input [31:0] result98,
	input [31:0] result99,
	input [31:0] result100,
	input [31:0] result101,
	input [31:0] result102,
	input [31:0] result103,
	input [31:0] result104,
	input [31:0] result105,
	input [31:0] result106,
	input [31:0] result107,
	input [31:0] result108,
	input [31:0] result109,
	input [31:0] result110,
	input [31:0] result111,
	input [31:0] result112,
	input [31:0] result113,
	input [31:0] result114,
	input [31:0] result115,
	input [31:0] result116,
	input [31:0] result117,
	input [31:0] result118,
	input [31:0] result119,
	input [31:0] result120,
	input [31:0] result121,
	input [31:0] result122,
	input [31:0] result123,
	input [31:0] result124,
	input [31:0] result125,
	input [31:0] result126,
	input [31:0] result127,
	input [31:0] result128,
	input [31:0] result129,
	input [31:0] result130,
	input [31:0] result131,
	input [31:0] result132,
	input [31:0] result133,
	input [31:0] result134,
	input [31:0] result135,
	input [31:0] result136,
	input [31:0] result137,
	input [31:0] result138,
	input [31:0] result139,
	input [31:0] result140,
	input [31:0] result141,
	input [31:0] result142,
	input [31:0] result143,
	input [31:0] result144,
	input [31:0] result145,
	input [31:0] result146,
	input [31:0] result147,
	input [31:0] result148,
	input [31:0] result149,
	input [31:0] result150,
	input [31:0] result151,
	input [31:0] result152,
	input [31:0] result153,
	input [31:0] result154,
	input [31:0] result155,
	input [31:0] result156,
	input [31:0] result157,
	input [31:0] result158,
	input [31:0] result159,
	input [31:0] result160,
	input [31:0] result161,
	input [31:0] result162,
	input [31:0] result163,
	input [31:0] result164,
	input [31:0] result165,
	input [31:0] result166,
	input [31:0] result167,
	input [31:0] result168,
	input [31:0] result169,
	input [31:0] result170,
	input [31:0] result171,
	input [31:0] result172,
	input [31:0] result173,
	input [31:0] result174,
	input [31:0] result175,
	input [31:0] result176,
	input [31:0] result177,
	input [31:0] result178,
	input [31:0] result179,
	input [31:0] result180,
	input [31:0] result181,
	input [31:0] result182,
	input [31:0] result183,
	input [31:0] result184,
	input [31:0] result185,
	input [31:0] result186,
	input [31:0] result187,
	input [31:0] result188,
	input [31:0] result189,
	input [31:0] result190,
	input [31:0] result191,
	input [31:0] result192,
	input [31:0] result193,
	input [31:0] result194,
	input [31:0] result195,
	input [31:0] result196,
	input [31:0] result197,
	input [31:0] result198,
	input [31:0] result199,
	input [31:0] result200,
	input [31:0] result201,
	input [31:0] result202,
	input [31:0] result203,
	input [31:0] result204,
	input [31:0] result205,
	input [31:0] result206,
	input [31:0] result207,
	input [31:0] result208,
	input [31:0] result209,
	input [31:0] result210,
	input [31:0] result211,
	input [31:0] result212,
	input [31:0] result213,
	input [31:0] result214,
	input [31:0] result215,
	input [31:0] result216,
	input [31:0] result217,
	input [31:0] result218,
	input [31:0] result219,
	input [31:0] result220,
	input [31:0] result221,
	input [31:0] result222,
	input [31:0] result223,
	input [31:0] result224,
	input [31:0] result225,
	input [31:0] result226,
	input [31:0] result227,
	input [31:0] result228,
	input [31:0] result229,
	input [31:0] result230,
	input [31:0] result231,
	input [31:0] result232,
	input [31:0] result233,
	input [31:0] result234,
	input [31:0] result235,
	input [31:0] result236,
	input [31:0] result237,
	input [31:0] result238,
	input [31:0] result239,
	input [31:0] result240,
	input [31:0] result241,
	input [31:0] result242,
	input [31:0] result243,
	input [31:0] result244,
	input [31:0] result245,
	input [31:0] result246,
	input [31:0] result247,
	input [31:0] result248,
	input [31:0] result249,
	input [31:0] result250,
	input [31:0] result251,
	input [31:0] result252,
	input [31:0] result253,
	input [31:0] result254,
	input [31:0] result255
);

	wire [7:0] counter;
	wire pim_status_read;
	wire busy, valid;

	wire weight_in_en, weight_out_en, weight_out_en_pim;
	wire [1:0] weight_sel;
	reg [8:0] WL_address;
	wire [8:0] WL_address_tmp;
	wire [31:0] weight_in_data;
	wire [255:0] cam_data;
	wire [255:0] cim_data;

	wire activation_in_en, activation_out_en, activation_out_en_pim;
	wire [1:0] activation_sel;
	wire [31:0] actvation_in_data;
	wire [287:0] activation_out_data;

	wire result_in_en, result_out_en, result_buffer_busy;
	wire [8191:0] result_in;
	wire [31:0] result_out;

	
	pim_controller controller(
		.i_clk						(i_clk), 
		.i_rst						(i_rst),
		.i_address					(i_address),

		.o_weight_in_en				(weight_in_en),	
		.o_weight_out_en			(weight_out_en),
		.o_weight_sel				(weight_sel),
		.o_WL_address				(WL_address_tmp),

		.o_activation_in_en			(activation_in_en),
		.o_activation_out_en		(activation_out_en),
		.o_activation_sel			(activation_sel),

		.o_result_buffer_busy		(result_buffer_busy),
		.o_result_in_en				(result_in_en),
		.o_result_out_en			(result_out_en),

		.o_counter					(counter),
		.o_busy						(busy),
		.o_valid					(valid),
		.o_pim_status_read					(pim_status_read)
	);

	weight_buffer WB (
		.i_clk						(i_clk),
		.i_rst						(i_rst),
		.i_weight_in_en				(weight_in_en),			
		.i_weight_out_en			(weight_out_en),
		.i_counter					(counter[3:0]),
		.i_data						(weight_in_data),
		.o_weight_out_en			(weight_out_en_pim),
		.o_cam_data					(cam_data),
		.o_cim_data					(cim_data)
	);

	activation_buffer AB (
		.i_clk						(i_clk),
		.i_rst						(i_rst),
		.i_activation_in_en			(activation_in_en),		
		.i_activation_out_en		(activation_out_en),
		.i_counter					(counter),
		.i_data						(actvation_in_data),
		.o_activation_out_en		(activation_out_en_pim),
		.o_data						(activation_out_data)
	);

	result_buffer RB(
		.i_clk						(i_clk),
		.i_rst						(i_rst),
		.i_result_buffer_busy		(result_buffer_busy),
		.i_result_in_en				(result_in_en),
		.i_result_out_en			(result_out_en),
		.i_counter					(counter),
		.i_data0					(result0),
		.i_data1					(result1),
		.i_data2					(result2),
		.i_data3					(result3),
		.i_data4					(result4),
		.i_data5					(result5),
		.i_data6					(result6),
		.i_data7					(result7),
		.i_data8					(result8),
		.i_data9					(result9),
		.i_data10					(result10),
		.i_data11					(result11),
		.i_data12					(result12),
		.i_data13					(result13),
		.i_data14					(result14),
		.i_data15					(result15),
		.i_data16					(result16),
		.i_data17					(result17),
		.i_data18					(result18),
		.i_data19					(result19),
		.i_data20					(result20),
		.i_data21					(result21),
		.i_data22					(result22),
		.i_data23					(result23),
		.i_data24					(result24),
		.i_data25					(result25),
		.i_data26					(result26),
		.i_data27					(result27),
		.i_data28					(result28),
		.i_data29					(result29),
		.i_data30					(result30),
		.i_data31					(result31),
		.i_data32					(result32),
		.i_data33					(result33),
		.i_data34					(result34),
		.i_data35					(result35),
		.i_data36					(result36),
		.i_data37					(result37),
		.i_data38					(result38),
		.i_data39					(result39),
		.i_data40					(result40),
		.i_data41					(result41),
		.i_data42					(result42),
		.i_data43					(result43),
		.i_data44					(result44),
		.i_data45					(result45),
		.i_data46					(result46),
		.i_data47					(result47),
		.i_data48					(result48),
		.i_data49					(result49),
		.i_data50					(result50),
		.i_data51					(result51),
		.i_data52					(result52),
		.i_data53					(result53),
		.i_data54					(result54),
		.i_data55					(result55),
		.i_data56					(result56),
		.i_data57					(result57),
		.i_data58					(result58),
		.i_data59					(result59),
		.i_data60					(result60),
		.i_data61					(result61),
		.i_data62					(result62),
		.i_data63					(result63),
		.i_data64					(result64),
		.i_data65					(result65),
		.i_data66					(result66),
		.i_data67					(result67),
		.i_data68					(result68),
		.i_data69					(result69),
		.i_data70					(result70),
		.i_data71					(result71),
		.i_data72					(result72),
		.i_data73					(result73),
		.i_data74					(result74),
		.i_data75					(result75),
		.i_data76					(result76),
		.i_data77					(result77),
		.i_data78					(result78),
		.i_data79					(result79),
		.i_data80					(result80),
		.i_data81					(result81),
		.i_data82					(result82),
		.i_data83					(result83),
		.i_data84					(result84),
		.i_data85					(result85),
		.i_data86					(result86),
		.i_data87					(result87),
		.i_data88					(result88),
		.i_data89					(result89),
		.i_data90					(result90),
		.i_data91					(result91),
		.i_data92					(result92),
		.i_data93					(result93),
		.i_data94					(result94),
		.i_data95					(result95),
		.i_data96					(result96),
		.i_data97					(result97),
		.i_data98					(result98),
		.i_data99					(result99),
		.i_data100					(result100),		
		.i_data101					(result101),
		.i_data102					(result102),
		.i_data103					(result103),
		.i_data104					(result104),
		.i_data105					(result105),
		.i_data106					(result106),
		.i_data107					(result107),
		.i_data108					(result108),
		.i_data109					(result109),
		.i_data110					(result110),
		.i_data111					(result111),
		.i_data112					(result112),
		.i_data113					(result113),
		.i_data114					(result114),
		.i_data115					(result115),
		.i_data116					(result116),
		.i_data117					(result117),
		.i_data118					(result118),
		.i_data119					(result119),
		.i_data120					(result120),
		.i_data121					(result121),
		.i_data122					(result122),
		.i_data123					(result123),
		.i_data124					(result124),
		.i_data125					(result125),
		.i_data126					(result126),
		.i_data127					(result127),
		.i_data128					(result128),
		.i_data129					(result129),
		.i_data130					(result130),
		.i_data131					(result131),
		.i_data132					(result132),
		.i_data133					(result133),
		.i_data134					(result134),
		.i_data135					(result135),
		.i_data136					(result136),
		.i_data137					(result137),
		.i_data138					(result138),
		.i_data139					(result139),
		.i_data140					(result140),
		.i_data141					(result141),
		.i_data142					(result142),
		.i_data143					(result143),
		.i_data144					(result144),
		.i_data145					(result145),
		.i_data146					(result146),
		.i_data147					(result147),
		.i_data148					(result148),
		.i_data149					(result149),
		.i_data150					(result150),
		.i_data151					(result151),
		.i_data152					(result152),
		.i_data153					(result153),
		.i_data154					(result154),
		.i_data155					(result155),
		.i_data156					(result156),
		.i_data157					(result157),
		.i_data158					(result158),
		.i_data159					(result159),
		.i_data160					(result160),
		.i_data161					(result161),
		.i_data162					(result162),
		.i_data163					(result163),
		.i_data164					(result164),
		.i_data165					(result165),
		.i_data166					(result166),
		.i_data167					(result167),
		.i_data168					(result168),
		.i_data169					(result169),
		.i_data170					(result170),
		.i_data171					(result171),
		.i_data172					(result172),
		.i_data173					(result173),
		.i_data174					(result174),
		.i_data175					(result175),
		.i_data176					(result176),
		.i_data177					(result177),
		.i_data178					(result178),
		.i_data179					(result179),
		.i_data180					(result180),
		.i_data181					(result181),
		.i_data182					(result182),
		.i_data183					(result183),
		.i_data184					(result184),
		.i_data185					(result185),
		.i_data186					(result186),
		.i_data187					(result187),
		.i_data188					(result188),
		.i_data189					(result189),
		.i_data190					(result190),
		.i_data191					(result191),
		.i_data192					(result192),
		.i_data193					(result193),
		.i_data194					(result194),
		.i_data195					(result195),
		.i_data196					(result196),
		.i_data197					(result197),
		.i_data198					(result198),
		.i_data199					(result199),
		.i_data200					(result200),
		.i_data201					(result201),
		.i_data202					(result202),
		.i_data203					(result203),
		.i_data204					(result204),
		.i_data205					(result205),
		.i_data206					(result206),
		.i_data207					(result207),
		.i_data208					(result208),
		.i_data209					(result209),
		.i_data210					(result210),
		.i_data211					(result211),
		.i_data212					(result212),
		.i_data213					(result213),
		.i_data214					(result214),
		.i_data215					(result215),
		.i_data216					(result216),
		.i_data217					(result217),
		.i_data218					(result218),
		.i_data219					(result219),
		.i_data220					(result220),
		.i_data221					(result221),
		.i_data222					(result222),
		.i_data223					(result223),
		.i_data224					(result224),
		.i_data225					(result225),
		.i_data226					(result226),
		.i_data227					(result227),
		.i_data228					(result228),
		.i_data229					(result229),
		.i_data230					(result230),
		.i_data231					(result231),
		.i_data232					(result232),
		.i_data233					(result233),
		.i_data234					(result234),
		.i_data235					(result235),
		.i_data236					(result236),
		.i_data237					(result237),
		.i_data238					(result238),
		.i_data239					(result239),
		.i_data240					(result240),
		.i_data241					(result241),
		.i_data242					(result242),
		.i_data243					(result243),
		.i_data244					(result244),
		.i_data245					(result245),
		.i_data246					(result246),
		.i_data247					(result247),
		.i_data248					(result248),
		.i_data249					(result249),
		.i_data250					(result250),
		.i_data251					(result251),
		.i_data252					(result252),
		.i_data253					(result253),
		.i_data254					(result254),
		.i_data255					(result255),
		.o_data						(result_out)
	);

	// dmux  #(
	// 	.width			(256)
	// ) cam_weight_sel (
	// 	.i_in			(cam_data),
	// 	.i_sel			(weight_sel),
	// 	.o_out0			(o_cam_data0),
	// 	.o_out1			(o_cam_data1),
	// 	.o_out2			(o_cam_data2),
	// 	.o_out3			(o_cam_data3)
	// );

	// dmux  #(
	// 	.width			(256)
	// ) cim_weight_sel (
	// 	.i_in			(cim_data),
	// 	.i_sel			(weight_sel),
	// 	.o_out0			(o_cim_data0),
	// 	.o_out1			(o_cim_data1),
	// 	.o_out2			(o_cim_data2),
	// 	.o_out3			(o_cim_data3)
	// );

	// dmux  #(
	// 	.width			(1)
	// ) weight_out_sel (
	// 	.i_in			(weight_out_en_pim),
	// 	.i_sel			(weight_sel),
	// 	.o_out0			(o_weight_out_en0),
	// 	.o_out1			(o_weight_out_en1),
	// 	.o_out2			(o_weight_out_en2),
	// 	.o_out3			(o_weight_out_en3)
	// );

	// dmux  #(
	// 	.width			(9)
	// ) WL_address_sel (
	// 	.i_in			(WL_address),
	// 	.i_sel			(weight_sel),
	// 	.o_out0			(o_WL_address0),
	// 	.o_out1			(o_WL_address1),
	// 	.o_out2			(o_WL_address2),
	// 	.o_out3			(o_WL_address3)
	// );

	// dmux  #(
	// 	.width			(1)
	// ) activation_out_sel (
	// 	.i_in			(activation_out_en_pim),
	// 	.i_sel			(activation_sel),
	// 	.o_out0			(o_activation_out_en0),
	// 	.o_out1			(o_activation_out_en1),
	// 	.o_out2			(o_activation_out_en2),
	// 	.o_out3			(o_activation_out_en3)
	// );

	// dmux  #(
	// 	.width			(288)
	// ) activation_out_data_sel (
	// 	.i_in			(activation_out_data),
	// 	.i_sel			(activation_sel),
	// 	.o_out0			(o_activation_out_data0),
	// 	.o_out1			(o_activation_out_data1),
	// 	.o_out2			(o_activation_out_data2),
	// 	.o_out3			(o_activation_out_data3)
	// );

	// mux #(
	// 	.width			(8192)
	// ) result_in_sel (
	// 	.i_in0			(i_result_in0),
	// 	.i_in1			(i_result_in1),
	// 	.i_in2			(i_result_in2),
	// 	.i_in3			(i_result_in3),
	// 	.i_sel			(activation_sel),
	// 	.o_out			(result_in)
	// );

	assign weight_in_data = weight_in_en ? i_data : 32'b0;
	assign actvation_in_data = activation_in_en ? i_data : 32'b0;

	// assign WL_address = weight_out_en ? WL_address_tmp : 9'd288;
	always @(posedge i_clk) begin
		if (i_rst) begin
			WL_address <= 0;
		end else begin
			if (weight_out_en) begin
				WL_address <= WL_address_tmp;
			end
		end
	end

	assign o_data = pim_status_read ? {30'b0, valid, busy} : result_out;

endmodule