module WL_driver (
	input i_pim_weight_in_en,
	input [8:0] i_WL_address,
	output reg [287:0] o_WL
);

	always @(*) begin
		if (i_pim_weight_in_en) begin
			case (i_WL_address) 
				9'd0  : begin o_WL[  0] = 1; o_WL[287:  1] = 0; end
				9'd1  : begin o_WL[  1] = 1; o_WL[287:  2] = 0; o_WL[0] = 0; end
				9'd2  : begin o_WL[  2] = 1; o_WL[287:  3] = 0; o_WL[  1:0] = 0; end
				9'd3  : begin o_WL[  3] = 1; o_WL[287:  4] = 0; o_WL[  2:0] = 0; end
				9'd4  : begin o_WL[  4] = 1; o_WL[287:  5] = 0; o_WL[  3:0] = 0; end
				9'd5  : begin o_WL[  5] = 1; o_WL[287:  6] = 0; o_WL[  4:0] = 0; end
				9'd6  : begin o_WL[  6] = 1; o_WL[287:  7] = 0; o_WL[  5:0] = 0; end
				9'd7  : begin o_WL[  7] = 1; o_WL[287:  8] = 0; o_WL[  6:0] = 0; end
				9'd8  : begin o_WL[  8] = 1; o_WL[287:  9] = 0; o_WL[  7:0] = 0; end
				9'd9  : begin o_WL[  9] = 1; o_WL[287: 10] = 0; o_WL[  8:0] = 0; end
				9'd10 : begin o_WL[ 10] = 1; o_WL[287: 11] = 0; o_WL[  9:0] = 0; end
				9'd11 : begin o_WL[ 11] = 1; o_WL[287: 12] = 0; o_WL[ 10:0] = 0; end
				9'd12 : begin o_WL[ 12] = 1; o_WL[287: 13] = 0; o_WL[ 11:0] = 0; end
				9'd13 : begin o_WL[ 13] = 1; o_WL[287: 14] = 0; o_WL[ 12:0] = 0; end
				9'd14 : begin o_WL[ 14] = 1; o_WL[287: 15] = 0; o_WL[ 13:0] = 0; end
				9'd15 : begin o_WL[ 15] = 1; o_WL[287: 16] = 0; o_WL[ 14:0] = 0; end
				9'd16 : begin o_WL[ 16] = 1; o_WL[287: 17] = 0; o_WL[ 15:0] = 0; end
				9'd17 : begin o_WL[ 17] = 1; o_WL[287: 18] = 0; o_WL[ 16:0] = 0; end
				9'd18 : begin o_WL[ 18] = 1; o_WL[287: 19] = 0; o_WL[ 17:0] = 0; end
				9'd19 : begin o_WL[ 19] = 1; o_WL[287: 20] = 0; o_WL[ 18:0] = 0; end
				9'd20 : begin o_WL[ 20] = 1; o_WL[287: 21] = 0; o_WL[ 19:0] = 0; end
				9'd21 : begin o_WL[ 21] = 1; o_WL[287: 22] = 0; o_WL[ 20:0] = 0; end
				9'd22 : begin o_WL[ 22] = 1; o_WL[287: 23] = 0; o_WL[ 21:0] = 0; end
				9'd23 : begin o_WL[ 23] = 1; o_WL[287: 24] = 0; o_WL[ 22:0] = 0; end
				9'd24 : begin o_WL[ 24] = 1; o_WL[287: 25] = 0; o_WL[ 23:0] = 0; end
				9'd25 : begin o_WL[ 25] = 1; o_WL[287: 26] = 0; o_WL[ 24:0] = 0; end
				9'd26 : begin o_WL[ 26] = 1; o_WL[287: 27] = 0; o_WL[ 25:0] = 0; end
				9'd27 : begin o_WL[ 27] = 1; o_WL[287: 28] = 0; o_WL[ 26:0] = 0; end
				9'd28 : begin o_WL[ 28] = 1; o_WL[287: 29] = 0; o_WL[ 27:0] = 0; end
				9'd29 : begin o_WL[ 29] = 1; o_WL[287: 30] = 0; o_WL[ 28:0] = 0; end
				9'd30 : begin o_WL[ 30] = 1; o_WL[287: 31] = 0; o_WL[ 29:0] = 0; end
				9'd31 : begin o_WL[ 31] = 1; o_WL[287: 32] = 0; o_WL[ 30:0] = 0; end
				9'd32 : begin o_WL[ 32] = 1; o_WL[287: 33] = 0; o_WL[ 31:0] = 0; end
				9'd33 : begin o_WL[ 33] = 1; o_WL[287: 34] = 0; o_WL[ 32:0] = 0; end
				9'd34 : begin o_WL[ 34] = 1; o_WL[287: 35] = 0; o_WL[ 33:0] = 0; end
				9'd35 : begin o_WL[ 35] = 1; o_WL[287: 36] = 0; o_WL[ 34:0] = 0; end
				9'd36 : begin o_WL[ 36] = 1; o_WL[287: 37] = 0; o_WL[ 35:0] = 0; end
				9'd37 : begin o_WL[ 37] = 1; o_WL[287: 38] = 0; o_WL[ 36:0] = 0; end
				9'd38 : begin o_WL[ 38] = 1; o_WL[287: 39] = 0; o_WL[ 37:0] = 0; end
				9'd39 : begin o_WL[ 39] = 1; o_WL[287: 40] = 0; o_WL[ 38:0] = 0; end
				9'd40 : begin o_WL[ 40] = 1; o_WL[287: 41] = 0; o_WL[ 39:0] = 0; end
				9'd41 : begin o_WL[ 41] = 1; o_WL[287: 42] = 0; o_WL[ 40:0] = 0; end
				9'd42 : begin o_WL[ 42] = 1; o_WL[287: 43] = 0; o_WL[ 41:0] = 0; end
				9'd43 : begin o_WL[ 43] = 1; o_WL[287: 44] = 0; o_WL[ 42:0] = 0; end
				9'd44 : begin o_WL[ 44] = 1; o_WL[287: 45] = 0; o_WL[ 43:0] = 0; end
				9'd45 : begin o_WL[ 45] = 1; o_WL[287: 46] = 0; o_WL[ 44:0] = 0; end
				9'd46 : begin o_WL[ 46] = 1; o_WL[287: 47] = 0; o_WL[ 45:0] = 0; end
				9'd47 : begin o_WL[ 47] = 1; o_WL[287: 48] = 0; o_WL[ 46:0] = 0; end
				9'd48 : begin o_WL[ 48] = 1; o_WL[287: 49] = 0; o_WL[ 47:0] = 0; end
				9'd49 : begin o_WL[ 49] = 1; o_WL[287: 50] = 0; o_WL[ 48:0] = 0; end
				9'd50 : begin o_WL[ 50] = 1; o_WL[287: 51] = 0; o_WL[ 49:0] = 0; end
				9'd51 : begin o_WL[ 51] = 1; o_WL[287: 52] = 0; o_WL[ 50:0] = 0; end
				9'd52 : begin o_WL[ 52] = 1; o_WL[287: 53] = 0; o_WL[ 51:0] = 0; end
				9'd53 : begin o_WL[ 53] = 1; o_WL[287: 54] = 0; o_WL[ 52:0] = 0; end
				9'd54 : begin o_WL[ 54] = 1; o_WL[287: 55] = 0; o_WL[ 53:0] = 0; end
				9'd55 : begin o_WL[ 55] = 1; o_WL[287: 56] = 0; o_WL[ 54:0] = 0; end
				9'd56 : begin o_WL[ 56] = 1; o_WL[287: 57] = 0; o_WL[ 55:0] = 0; end
				9'd57 : begin o_WL[ 57] = 1; o_WL[287: 58] = 0; o_WL[ 56:0] = 0; end
				9'd58 : begin o_WL[ 58] = 1; o_WL[287: 59] = 0; o_WL[ 57:0] = 0; end
				9'd59 : begin o_WL[ 59] = 1; o_WL[287: 60] = 0; o_WL[ 58:0] = 0; end
				9'd60 : begin o_WL[ 60] = 1; o_WL[287: 61] = 0; o_WL[ 59:0] = 0; end
				9'd61 : begin o_WL[ 61] = 1; o_WL[287: 62] = 0; o_WL[ 60:0] = 0; end
				9'd62 : begin o_WL[ 62] = 1; o_WL[287: 63] = 0; o_WL[ 61:0] = 0; end
				9'd63 : begin o_WL[ 63] = 1; o_WL[287: 64] = 0; o_WL[ 62:0] = 0; end
				9'd64 : begin o_WL[ 64] = 1; o_WL[287: 65] = 0; o_WL[ 63:0] = 0; end
				9'd65 : begin o_WL[ 65] = 1; o_WL[287: 66] = 0; o_WL[ 64:0] = 0; end
				9'd66 : begin o_WL[ 66] = 1; o_WL[287: 67] = 0; o_WL[ 65:0] = 0; end
				9'd67 : begin o_WL[ 67] = 1; o_WL[287: 68] = 0; o_WL[ 66:0] = 0; end
				9'd68 : begin o_WL[ 68] = 1; o_WL[287: 69] = 0; o_WL[ 67:0] = 0; end
				9'd69 : begin o_WL[ 69] = 1; o_WL[287: 70] = 0; o_WL[ 68:0] = 0; end
				9'd70 : begin o_WL[ 70] = 1; o_WL[287: 71] = 0; o_WL[ 69:0] = 0; end
				9'd71 : begin o_WL[ 71] = 1; o_WL[287: 72] = 0; o_WL[ 70:0] = 0; end
				9'd72 : begin o_WL[ 72] = 1; o_WL[287: 73] = 0; o_WL[ 71:0] = 0; end
				9'd73 : begin o_WL[ 73] = 1; o_WL[287: 74] = 0; o_WL[ 72:0] = 0; end
				9'd74 : begin o_WL[ 74] = 1; o_WL[287: 75] = 0; o_WL[ 73:0] = 0; end
				9'd75 : begin o_WL[ 75] = 1; o_WL[287: 76] = 0; o_WL[ 74:0] = 0; end
				9'd76 : begin o_WL[ 76] = 1; o_WL[287: 77] = 0; o_WL[ 75:0] = 0; end
				9'd77 : begin o_WL[ 77] = 1; o_WL[287: 78] = 0; o_WL[ 76:0] = 0; end
				9'd78 : begin o_WL[ 78] = 1; o_WL[287: 79] = 0; o_WL[ 77:0] = 0; end
				9'd79 : begin o_WL[ 79] = 1; o_WL[287: 80] = 0; o_WL[ 78:0] = 0; end
				9'd80 : begin o_WL[ 80] = 1; o_WL[287: 81] = 0; o_WL[ 79:0] = 0; end
				9'd81 : begin o_WL[ 81] = 1; o_WL[287: 82] = 0; o_WL[ 80:0] = 0; end
				9'd82 : begin o_WL[ 82] = 1; o_WL[287: 83] = 0; o_WL[ 81:0] = 0; end
				9'd83 : begin o_WL[ 83] = 1; o_WL[287: 84] = 0; o_WL[ 82:0] = 0; end
				9'd84 : begin o_WL[ 84] = 1; o_WL[287: 85] = 0; o_WL[ 83:0] = 0; end
				9'd85 : begin o_WL[ 85] = 1; o_WL[287: 86] = 0; o_WL[ 84:0] = 0; end
				9'd86 : begin o_WL[ 86] = 1; o_WL[287: 87] = 0; o_WL[ 85:0] = 0; end
				9'd87 : begin o_WL[ 87] = 1; o_WL[287: 88] = 0; o_WL[ 86:0] = 0; end
				9'd88 : begin o_WL[ 88] = 1; o_WL[287: 89] = 0; o_WL[ 87:0] = 0; end
				9'd89 : begin o_WL[ 89] = 1; o_WL[287: 90] = 0; o_WL[ 88:0] = 0; end
				9'd90 : begin o_WL[ 90] = 1; o_WL[287: 91] = 0; o_WL[ 89:0] = 0; end
				9'd91 : begin o_WL[ 91] = 1; o_WL[287: 92] = 0; o_WL[ 90:0] = 0; end
				9'd92 : begin o_WL[ 92] = 1; o_WL[287: 93] = 0; o_WL[ 91:0] = 0; end
				9'd93 : begin o_WL[ 93] = 1; o_WL[287: 94] = 0; o_WL[ 92:0] = 0; end
				9'd94 : begin o_WL[ 94] = 1; o_WL[287: 95] = 0; o_WL[ 93:0] = 0; end
				9'd95 : begin o_WL[ 95] = 1; o_WL[287: 96] = 0; o_WL[ 94:0] = 0; end
				9'd96 : begin o_WL[ 96] = 1; o_WL[287: 97] = 0; o_WL[ 95:0] = 0; end
				9'd97 : begin o_WL[ 97] = 1; o_WL[287: 98] = 0; o_WL[ 96:0] = 0; end
				9'd98 : begin o_WL[ 98] = 1; o_WL[287: 99] = 0; o_WL[ 97:0] = 0; end
				9'd99 : begin o_WL[ 99] = 1; o_WL[287:100] = 0; o_WL[ 98:0] = 0; end
				9'd100: begin o_WL[100] = 1; o_WL[287:101] = 0; o_WL[ 99:0] = 0; end
				9'd101: begin o_WL[101] = 1; o_WL[287:102] = 0; o_WL[100:0] = 0; end
				9'd102: begin o_WL[102] = 1; o_WL[287:103] = 0; o_WL[101:0] = 0; end
				9'd103: begin o_WL[103] = 1; o_WL[287:104] = 0; o_WL[102:0] = 0; end
				9'd104: begin o_WL[104] = 1; o_WL[287:105] = 0; o_WL[103:0] = 0; end
				9'd105: begin o_WL[105] = 1; o_WL[287:106] = 0; o_WL[104:0] = 0; end
				9'd106: begin o_WL[106] = 1; o_WL[287:107] = 0; o_WL[105:0] = 0; end
				9'd107: begin o_WL[107] = 1; o_WL[287:108] = 0; o_WL[106:0] = 0; end
				9'd108: begin o_WL[108] = 1; o_WL[287:109] = 0; o_WL[107:0] = 0; end
				9'd109: begin o_WL[109] = 1; o_WL[287:110] = 0; o_WL[108:0] = 0; end
				9'd110: begin o_WL[110] = 1; o_WL[287:111] = 0; o_WL[109:0] = 0; end
				9'd111: begin o_WL[111] = 1; o_WL[287:112] = 0; o_WL[110:0] = 0; end
				9'd112: begin o_WL[112] = 1; o_WL[287:113] = 0; o_WL[111:0] = 0; end
				9'd113: begin o_WL[113] = 1; o_WL[287:114] = 0; o_WL[112:0] = 0; end
				9'd114: begin o_WL[114] = 1; o_WL[287:115] = 0; o_WL[113:0] = 0; end
				9'd115: begin o_WL[115] = 1; o_WL[287:116] = 0; o_WL[114:0] = 0; end
				9'd116: begin o_WL[116] = 1; o_WL[287:117] = 0; o_WL[115:0] = 0; end
				9'd117: begin o_WL[117] = 1; o_WL[287:118] = 0; o_WL[116:0] = 0; end
				9'd118: begin o_WL[118] = 1; o_WL[287:119] = 0; o_WL[117:0] = 0; end
				9'd119: begin o_WL[119] = 1; o_WL[287:120] = 0; o_WL[118:0] = 0; end
				9'd120: begin o_WL[120] = 1; o_WL[287:121] = 0; o_WL[119:0] = 0; end
				9'd121: begin o_WL[121] = 1; o_WL[287:122] = 0; o_WL[120:0] = 0; end
				9'd122: begin o_WL[122] = 1; o_WL[287:123] = 0; o_WL[121:0] = 0; end
				9'd123: begin o_WL[123] = 1; o_WL[287:124] = 0; o_WL[122:0] = 0; end
				9'd124: begin o_WL[124] = 1; o_WL[287:125] = 0; o_WL[123:0] = 0; end
				9'd125: begin o_WL[125] = 1; o_WL[287:126] = 0; o_WL[124:0] = 0; end
				9'd126: begin o_WL[126] = 1; o_WL[287:127] = 0; o_WL[125:0] = 0; end
				9'd127: begin o_WL[127] = 1; o_WL[287:128] = 0; o_WL[126:0] = 0; end
				9'd128: begin o_WL[128] = 1; o_WL[287:129] = 0; o_WL[127:0] = 0; end
				9'd129: begin o_WL[129] = 1; o_WL[287:130] = 0; o_WL[128:0] = 0; end
				9'd130: begin o_WL[130] = 1; o_WL[287:131] = 0; o_WL[129:0] = 0; end
				9'd131: begin o_WL[131] = 1; o_WL[287:132] = 0; o_WL[130:0] = 0; end
				9'd132: begin o_WL[132] = 1; o_WL[287:133] = 0; o_WL[131:0] = 0; end
				9'd133: begin o_WL[133] = 1; o_WL[287:134] = 0; o_WL[132:0] = 0; end
				9'd134: begin o_WL[134] = 1; o_WL[287:135] = 0; o_WL[133:0] = 0; end
				9'd135: begin o_WL[135] = 1; o_WL[287:136] = 0; o_WL[134:0] = 0; end
				9'd136: begin o_WL[136] = 1; o_WL[287:137] = 0; o_WL[135:0] = 0; end
				9'd137: begin o_WL[137] = 1; o_WL[287:138] = 0; o_WL[136:0] = 0; end
				9'd138: begin o_WL[138] = 1; o_WL[287:139] = 0; o_WL[137:0] = 0; end
				9'd139: begin o_WL[139] = 1; o_WL[287:140] = 0; o_WL[138:0] = 0; end
				9'd140: begin o_WL[140] = 1; o_WL[287:141] = 0; o_WL[139:0] = 0; end
				9'd141: begin o_WL[141] = 1; o_WL[287:142] = 0; o_WL[140:0] = 0; end
				9'd142: begin o_WL[142] = 1; o_WL[287:143] = 0; o_WL[141:0] = 0; end
				9'd143: begin o_WL[143] = 1; o_WL[287:144] = 0; o_WL[142:0] = 0; end
				9'd144: begin o_WL[144] = 1; o_WL[287:145] = 0; o_WL[143:0] = 0; end
				9'd145: begin o_WL[145] = 1; o_WL[287:146] = 0; o_WL[144:0] = 0; end
				9'd146: begin o_WL[146] = 1; o_WL[287:147] = 0; o_WL[145:0] = 0; end
				9'd147: begin o_WL[147] = 1; o_WL[287:148] = 0; o_WL[146:0] = 0; end
				9'd148: begin o_WL[148] = 1; o_WL[287:149] = 0; o_WL[147:0] = 0; end
				9'd149: begin o_WL[149] = 1; o_WL[287:150] = 0; o_WL[148:0] = 0; end
				9'd150: begin o_WL[150] = 1; o_WL[287:151] = 0; o_WL[149:0] = 0; end
				9'd151: begin o_WL[151] = 1; o_WL[287:152] = 0; o_WL[150:0] = 0; end
				9'd152: begin o_WL[152] = 1; o_WL[287:153] = 0; o_WL[151:0] = 0; end
				9'd153: begin o_WL[153] = 1; o_WL[287:154] = 0; o_WL[152:0] = 0; end
				9'd154: begin o_WL[154] = 1; o_WL[287:155] = 0; o_WL[153:0] = 0; end
				9'd155: begin o_WL[155] = 1; o_WL[287:156] = 0; o_WL[154:0] = 0; end
				9'd156: begin o_WL[156] = 1; o_WL[287:157] = 0; o_WL[155:0] = 0; end
				9'd157: begin o_WL[157] = 1; o_WL[287:158] = 0; o_WL[156:0] = 0; end
				9'd158: begin o_WL[158] = 1; o_WL[287:159] = 0; o_WL[157:0] = 0; end
				9'd159: begin o_WL[159] = 1; o_WL[287:160] = 0; o_WL[158:0] = 0; end
				9'd160: begin o_WL[160] = 1; o_WL[287:161] = 0; o_WL[159:0] = 0; end
				9'd161: begin o_WL[161] = 1; o_WL[287:162] = 0; o_WL[160:0] = 0; end
				9'd162: begin o_WL[162] = 1; o_WL[287:163] = 0; o_WL[161:0] = 0; end
				9'd163: begin o_WL[163] = 1; o_WL[287:164] = 0; o_WL[162:0] = 0; end
				9'd164: begin o_WL[164] = 1; o_WL[287:165] = 0; o_WL[163:0] = 0; end
				9'd165: begin o_WL[165] = 1; o_WL[287:166] = 0; o_WL[164:0] = 0; end
				9'd166: begin o_WL[166] = 1; o_WL[287:167] = 0; o_WL[165:0] = 0; end
				9'd167: begin o_WL[167] = 1; o_WL[287:168] = 0; o_WL[166:0] = 0; end
				9'd168: begin o_WL[168] = 1; o_WL[287:169] = 0; o_WL[167:0] = 0; end
				9'd169: begin o_WL[169] = 1; o_WL[287:170] = 0; o_WL[168:0] = 0; end
				9'd170: begin o_WL[170] = 1; o_WL[287:171] = 0; o_WL[169:0] = 0; end
				9'd171: begin o_WL[171] = 1; o_WL[287:172] = 0; o_WL[170:0] = 0; end
				9'd172: begin o_WL[172] = 1; o_WL[287:173] = 0; o_WL[171:0] = 0; end
				9'd173: begin o_WL[173] = 1; o_WL[287:174] = 0; o_WL[172:0] = 0; end
				9'd174: begin o_WL[174] = 1; o_WL[287:175] = 0; o_WL[173:0] = 0; end
				9'd175: begin o_WL[175] = 1; o_WL[287:176] = 0; o_WL[174:0] = 0; end
				9'd176: begin o_WL[176] = 1; o_WL[287:177] = 0; o_WL[175:0] = 0; end
				9'd177: begin o_WL[177] = 1; o_WL[287:178] = 0; o_WL[176:0] = 0; end
				9'd178: begin o_WL[178] = 1; o_WL[287:179] = 0; o_WL[177:0] = 0; end
				9'd179: begin o_WL[179] = 1; o_WL[287:180] = 0; o_WL[178:0] = 0; end
				9'd180: begin o_WL[180] = 1; o_WL[287:181] = 0; o_WL[179:0] = 0; end
				9'd181: begin o_WL[181] = 1; o_WL[287:182] = 0; o_WL[180:0] = 0; end
				9'd182: begin o_WL[182] = 1; o_WL[287:183] = 0; o_WL[181:0] = 0; end
				9'd183: begin o_WL[183] = 1; o_WL[287:184] = 0; o_WL[182:0] = 0; end
				9'd184: begin o_WL[184] = 1; o_WL[287:185] = 0; o_WL[183:0] = 0; end
				9'd185: begin o_WL[185] = 1; o_WL[287:186] = 0; o_WL[184:0] = 0; end
				9'd186: begin o_WL[186] = 1; o_WL[287:187] = 0; o_WL[185:0] = 0; end
				9'd187: begin o_WL[187] = 1; o_WL[287:188] = 0; o_WL[186:0] = 0; end
				9'd188: begin o_WL[188] = 1; o_WL[287:189] = 0; o_WL[187:0] = 0; end
				9'd189: begin o_WL[189] = 1; o_WL[287:190] = 0; o_WL[188:0] = 0; end
				9'd190: begin o_WL[190] = 1; o_WL[287:191] = 0; o_WL[189:0] = 0; end
				9'd191: begin o_WL[191] = 1; o_WL[287:192] = 0; o_WL[190:0] = 0; end
				9'd192: begin o_WL[192] = 1; o_WL[287:193] = 0; o_WL[191:0] = 0; end
				9'd193: begin o_WL[193] = 1; o_WL[287:194] = 0; o_WL[192:0] = 0; end
				9'd194: begin o_WL[194] = 1; o_WL[287:195] = 0; o_WL[193:0] = 0; end
				9'd195: begin o_WL[195] = 1; o_WL[287:196] = 0; o_WL[194:0] = 0; end
				9'd196: begin o_WL[196] = 1; o_WL[287:197] = 0; o_WL[195:0] = 0; end
				9'd197: begin o_WL[197] = 1; o_WL[287:198] = 0; o_WL[196:0] = 0; end
				9'd198: begin o_WL[198] = 1; o_WL[287:199] = 0; o_WL[197:0] = 0; end
				9'd199: begin o_WL[199] = 1; o_WL[287:200] = 0; o_WL[198:0] = 0; end
				9'd200: begin o_WL[200] = 1; o_WL[287:201] = 0; o_WL[199:0] = 0; end
				9'd201: begin o_WL[201] = 1; o_WL[287:202] = 0; o_WL[200:0] = 0; end
				9'd202: begin o_WL[202] = 1; o_WL[287:203] = 0; o_WL[201:0] = 0; end
				9'd203: begin o_WL[203] = 1; o_WL[287:204] = 0; o_WL[202:0] = 0; end
				9'd204: begin o_WL[204] = 1; o_WL[287:205] = 0; o_WL[203:0] = 0; end
				9'd205: begin o_WL[205] = 1; o_WL[287:206] = 0; o_WL[204:0] = 0; end
				9'd206: begin o_WL[206] = 1; o_WL[287:207] = 0; o_WL[205:0] = 0; end
				9'd207: begin o_WL[207] = 1; o_WL[287:208] = 0; o_WL[206:0] = 0; end
				9'd208: begin o_WL[208] = 1; o_WL[287:209] = 0; o_WL[207:0] = 0; end
				9'd209: begin o_WL[209] = 1; o_WL[287:210] = 0; o_WL[208:0] = 0; end
				9'd210: begin o_WL[210] = 1; o_WL[287:211] = 0; o_WL[209:0] = 0; end
				9'd211: begin o_WL[211] = 1; o_WL[287:212] = 0; o_WL[210:0] = 0; end
				9'd212: begin o_WL[212] = 1; o_WL[287:213] = 0; o_WL[211:0] = 0; end
				9'd213: begin o_WL[213] = 1; o_WL[287:214] = 0; o_WL[212:0] = 0; end
				9'd214: begin o_WL[214] = 1; o_WL[287:215] = 0; o_WL[213:0] = 0; end
				9'd215: begin o_WL[215] = 1; o_WL[287:216] = 0; o_WL[214:0] = 0; end
				9'd216: begin o_WL[216] = 1; o_WL[287:217] = 0; o_WL[215:0] = 0; end
				9'd217: begin o_WL[217] = 1; o_WL[287:218] = 0; o_WL[216:0] = 0; end
				9'd218: begin o_WL[218] = 1; o_WL[287:219] = 0; o_WL[217:0] = 0; end
				9'd219: begin o_WL[219] = 1; o_WL[287:220] = 0; o_WL[218:0] = 0; end
				9'd220: begin o_WL[220] = 1; o_WL[287:221] = 0; o_WL[219:0] = 0; end
				9'd221: begin o_WL[221] = 1; o_WL[287:222] = 0; o_WL[220:0] = 0; end
				9'd222: begin o_WL[222] = 1; o_WL[287:223] = 0; o_WL[221:0] = 0; end
				9'd223: begin o_WL[223] = 1; o_WL[287:224] = 0; o_WL[222:0] = 0; end
				9'd224: begin o_WL[224] = 1; o_WL[287:225] = 0; o_WL[223:0] = 0; end
				9'd225: begin o_WL[225] = 1; o_WL[287:226] = 0; o_WL[224:0] = 0; end
				9'd226: begin o_WL[226] = 1; o_WL[287:227] = 0; o_WL[225:0] = 0; end
				9'd227: begin o_WL[227] = 1; o_WL[287:228] = 0; o_WL[226:0] = 0; end
				9'd228: begin o_WL[228] = 1; o_WL[287:229] = 0; o_WL[227:0] = 0; end
				9'd229: begin o_WL[229] = 1; o_WL[287:230] = 0; o_WL[228:0] = 0; end
				9'd230: begin o_WL[230] = 1; o_WL[287:231] = 0; o_WL[229:0] = 0; end
				9'd231: begin o_WL[231] = 1; o_WL[287:232] = 0; o_WL[230:0] = 0; end
				9'd232: begin o_WL[232] = 1; o_WL[287:233] = 0; o_WL[231:0] = 0; end
				9'd233: begin o_WL[233] = 1; o_WL[287:234] = 0; o_WL[232:0] = 0; end
				9'd234: begin o_WL[234] = 1; o_WL[287:235] = 0; o_WL[233:0] = 0; end
				9'd235: begin o_WL[235] = 1; o_WL[287:236] = 0; o_WL[234:0] = 0; end
				9'd236: begin o_WL[236] = 1; o_WL[287:237] = 0; o_WL[235:0] = 0; end
				9'd237: begin o_WL[237] = 1; o_WL[287:238] = 0; o_WL[236:0] = 0; end
				9'd238: begin o_WL[238] = 1; o_WL[287:239] = 0; o_WL[237:0] = 0; end
				9'd239: begin o_WL[239] = 1; o_WL[287:240] = 0; o_WL[238:0] = 0; end
				9'd240: begin o_WL[240] = 1; o_WL[287:241] = 0; o_WL[239:0] = 0; end
				9'd241: begin o_WL[241] = 1; o_WL[287:242] = 0; o_WL[240:0] = 0; end
				9'd242: begin o_WL[242] = 1; o_WL[287:243] = 0; o_WL[241:0] = 0; end
				9'd243: begin o_WL[243] = 1; o_WL[287:244] = 0; o_WL[242:0] = 0; end
				9'd244: begin o_WL[244] = 1; o_WL[287:245] = 0; o_WL[243:0] = 0; end
				9'd245: begin o_WL[245] = 1; o_WL[287:246] = 0; o_WL[244:0] = 0; end
				9'd246: begin o_WL[246] = 1; o_WL[287:247] = 0; o_WL[245:0] = 0; end
				9'd247: begin o_WL[247] = 1; o_WL[287:248] = 0; o_WL[246:0] = 0; end
				9'd248: begin o_WL[248] = 1; o_WL[287:249] = 0; o_WL[247:0] = 0; end
				9'd249: begin o_WL[249] = 1; o_WL[287:250] = 0; o_WL[248:0] = 0; end
				9'd250: begin o_WL[250] = 1; o_WL[287:251] = 0; o_WL[249:0] = 0; end
				9'd251: begin o_WL[251] = 1; o_WL[287:252] = 0; o_WL[250:0] = 0; end
				9'd252: begin o_WL[252] = 1; o_WL[287:253] = 0; o_WL[251:0] = 0; end
				9'd253: begin o_WL[253] = 1; o_WL[287:254] = 0; o_WL[252:0] = 0; end
				9'd254: begin o_WL[254] = 1; o_WL[287:255] = 0; o_WL[253:0] = 0; end
				9'd255: begin o_WL[255] = 1; o_WL[287:256] = 0; o_WL[254:0] = 0; end
				9'd256: begin o_WL[256] = 1; o_WL[287:257] = 0; o_WL[255:0] = 0; end
				9'd257: begin o_WL[257] = 1; o_WL[287:258] = 0; o_WL[256:0] = 0; end
				9'd258: begin o_WL[258] = 1; o_WL[287:259] = 0; o_WL[257:0] = 0; end
				9'd259: begin o_WL[259] = 1; o_WL[287:260] = 0; o_WL[258:0] = 0; end
				9'd260: begin o_WL[260] = 1; o_WL[287:261] = 0; o_WL[259:0] = 0; end
				9'd261: begin o_WL[261] = 1; o_WL[287:262] = 0; o_WL[260:0] = 0; end
				9'd262: begin o_WL[262] = 1; o_WL[287:263] = 0; o_WL[261:0] = 0; end
				9'd263: begin o_WL[263] = 1; o_WL[287:264] = 0; o_WL[262:0] = 0; end
				9'd264: begin o_WL[264] = 1; o_WL[287:265] = 0; o_WL[263:0] = 0; end
				9'd265: begin o_WL[265] = 1; o_WL[287:266] = 0; o_WL[264:0] = 0; end
				9'd266: begin o_WL[266] = 1; o_WL[287:267] = 0; o_WL[265:0] = 0; end
				9'd267: begin o_WL[267] = 1; o_WL[287:268] = 0; o_WL[266:0] = 0; end
				9'd268: begin o_WL[268] = 1; o_WL[287:269] = 0; o_WL[267:0] = 0; end
				9'd269: begin o_WL[269] = 1; o_WL[287:270] = 0; o_WL[268:0] = 0; end
				9'd270: begin o_WL[270] = 1; o_WL[287:271] = 0; o_WL[269:0] = 0; end
				9'd271: begin o_WL[271] = 1; o_WL[287:272] = 0; o_WL[270:0] = 0; end
				9'd272: begin o_WL[272] = 1; o_WL[287:273] = 0; o_WL[271:0] = 0; end
				9'd273: begin o_WL[273] = 1; o_WL[287:274] = 0; o_WL[272:0] = 0; end
				9'd274: begin o_WL[274] = 1; o_WL[287:275] = 0; o_WL[273:0] = 0; end
				9'd275: begin o_WL[275] = 1; o_WL[287:276] = 0; o_WL[274:0] = 0; end
				9'd276: begin o_WL[276] = 1; o_WL[287:277] = 0; o_WL[275:0] = 0; end
				9'd277: begin o_WL[277] = 1; o_WL[287:278] = 0; o_WL[276:0] = 0; end
				9'd278: begin o_WL[278] = 1; o_WL[287:279] = 0; o_WL[277:0] = 0; end
				9'd279: begin o_WL[279] = 1; o_WL[287:280] = 0; o_WL[278:0] = 0; end
				9'd280: begin o_WL[280] = 1; o_WL[287:281] = 0; o_WL[279:0] = 0; end
				9'd281: begin o_WL[281] = 1; o_WL[287:282] = 0; o_WL[280:0] = 0; end
				9'd282: begin o_WL[282] = 1; o_WL[287:283] = 0; o_WL[281:0] = 0; end
				9'd283: begin o_WL[283] = 1; o_WL[287:284] = 0; o_WL[282:0] = 0; end
				9'd284: begin o_WL[284] = 1; o_WL[287:285] = 0; o_WL[283:0] = 0; end
				9'd285: begin o_WL[285] = 1; o_WL[287:286] = 0; o_WL[284:0] = 0; end
				9'd286: begin o_WL[286] = 1; o_WL[287] = 0; o_WL[285:0] = 0; end
				9'd287: begin o_WL[287] = 1;  o_WL[286:0] = 0; end 
				default: o_WL = 0;
			endcase	
		end 
	end


endmodule